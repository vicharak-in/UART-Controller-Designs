
//
// Verific Verilog Description of module UART_Controller
//

module UART_Controller (clk, rx, tx1, tx2, led_command, led_data, 
            jtag_inst1_CAPTURE, jtag_inst1_DRCK, jtag_inst1_RESET, jtag_inst1_RUNTEST, 
            jtag_inst1_SEL, jtag_inst1_SHIFT, jtag_inst1_TCK, jtag_inst1_TDI, 
            jtag_inst1_TMS, jtag_inst1_UPDATE, jtag_inst1_TDO);
    input clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input rx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output tx1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output tx2 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output led_command /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output led_data /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input jtag_inst1_CAPTURE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_DRCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RESET /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_RUNTEST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SEL /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_SHIFT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TCK /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TDI /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_TMS /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input jtag_inst1_UPDATE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output jtag_inst1_TDO /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    wire n257_2;
    wire n62_2;
    wire n61_2;
    wire n60_2;
    wire n59_2;
    wire n58_2;
    
    wire \data[0] , DV, \i[0] , \transmitter_select[0] , \data_length[0] , 
        \uart_rx/r_Clock_Count[0] , RX_DV, \uart_rx/r_RX_Byte[0] , \uart_rx/r_Bit_Index[0] , 
        \uart_rx/r_SM_Main[0] , \uart_rx/r_Clock_Count[1] , \uart_rx/r_Clock_Count[2] , 
        \uart_rx/r_Clock_Count[3] , \uart_rx/r_Clock_Count[4] , \uart_rx/r_Clock_Count[5] , 
        \uart_rx/r_Clock_Count[6] , \uart_rx/r_Clock_Count[7] , \uart_rx/r_RX_Byte[1] , 
        \uart_rx/r_RX_Byte[2] , \uart_rx/r_RX_Byte[3] , \uart_rx/r_RX_Byte[4] , 
        \uart_rx/r_RX_Byte[5] , \uart_rx/r_RX_Byte[6] , \uart_rx/r_RX_Byte[7] , 
        \uart_rx/r_Bit_Index[1] , \uart_rx/r_Bit_Index[2] , \uart_rx/r_SM_Main[1] , 
        \data[1] , \data[2] , \data[3] , \data[4] , \data[5] , \data[6] , 
        \data[7] , \i[1] , \i[2] , \i[3] , \i[4] , \i[5] , \transmitter_select[1] , 
        \data_length[1] , \data_length[2] , \data_length[3] , \data_length[4] , 
        \data_length[5] , \uart_tx1/r_Clock_Count[0] , \uart_tx1/r_Bit_Index[0] , 
        \uart_tx1/r_TX_Data[0] , \uart_tx1/r_SM_Main[0] , \uart_tx1/r_Clock_Count[1] , 
        \uart_tx1/r_Clock_Count[2] , \uart_tx1/r_Clock_Count[3] , \uart_tx1/r_Clock_Count[4] , 
        \uart_tx1/r_Clock_Count[5] , \uart_tx1/r_Clock_Count[6] , \uart_tx1/r_Bit_Index[1] , 
        \uart_tx1/r_Bit_Index[2] , \uart_tx1/r_TX_Data[1] , \uart_tx1/r_TX_Data[2] , 
        \uart_tx1/r_TX_Data[3] , \uart_tx1/r_TX_Data[4] , \uart_tx1/r_TX_Data[5] , 
        \uart_tx1/r_TX_Data[6] , \uart_tx1/r_TX_Data[7] , \uart_tx1/r_SM_Main[1] , 
        \uart_tx2/r_TX_Data[0] , \uart_tx2/r_TX_Data[1] , \uart_tx2/r_TX_Data[2] , 
        \uart_tx2/r_TX_Data[3] , \uart_tx2/r_TX_Data[4] , \uart_tx2/r_TX_Data[5] , 
        \uart_tx2/r_TX_Data[6] , \uart_tx2/r_TX_Data[7] , \edb_top_inst/n2270 , 
        \edb_top_inst/la0/la_run_trig , \edb_top_inst/la0/la_trig_pattern[0] , 
        \edb_top_inst/la0/la_run_trig_imdt , \edb_top_inst/la0/la_stop_trig , 
        \edb_top_inst/la0/la_capture_pattern[0] , \edb_top_inst/la0/la_trig_mask[0] , 
        \edb_top_inst/la0/la_num_trigger[0] , \edb_top_inst/la0/la_window_depth[0] , 
        \edb_top_inst/la0/la_soft_reset_in , \edb_top_inst/la0/address_counter[0] , 
        \edb_top_inst/la0/opcode[0] , \edb_top_inst/la0/bit_count[0] , \edb_top_inst/la0/word_count[0] , 
        \edb_top_inst/la0/data_out_shift_reg[0] , \edb_top_inst/la0/module_state[0] , 
        \edb_top_inst/la0/la_resetn_p1 , \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] , 
        \edb_top_inst/la0/la_resetn , \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] , \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] , 
        \edb_top_inst/la0/genblk2.la_capture_mask[0] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[0] , 
        \edb_top_inst/la0/cap_fifo_din_cu[1] , \edb_top_inst/la0/cap_fifo_din_cu[0] , 
        \edb_top_inst/la0/cap_fifo_din_tu[0] , \edb_top_inst/la0/internal_register_select[0] , 
        \edb_top_inst/la0/la_trig_pos[0] , \edb_top_inst/la0/la_trig_pattern[1] , 
        \edb_top_inst/la0/la_capture_pattern[1] , \edb_top_inst/la0/la_trig_mask[1] , 
        \edb_top_inst/la0/la_trig_mask[2] , \edb_top_inst/la0/la_trig_mask[3] , 
        \edb_top_inst/la0/la_trig_mask[4] , \edb_top_inst/la0/la_trig_mask[5] , 
        \edb_top_inst/la0/la_trig_mask[6] , \edb_top_inst/la0/la_trig_mask[7] , 
        \edb_top_inst/la0/la_trig_mask[8] , \edb_top_inst/la0/la_trig_mask[9] , 
        \edb_top_inst/la0/la_trig_mask[10] , \edb_top_inst/la0/la_trig_mask[11] , 
        \edb_top_inst/la0/la_trig_mask[12] , \edb_top_inst/la0/la_trig_mask[13] , 
        \edb_top_inst/la0/la_trig_mask[14] , \edb_top_inst/la0/la_trig_mask[15] , 
        \edb_top_inst/la0/la_trig_mask[16] , \edb_top_inst/la0/la_trig_mask[17] , 
        \edb_top_inst/la0/la_trig_mask[18] , \edb_top_inst/la0/la_trig_mask[19] , 
        \edb_top_inst/la0/la_trig_mask[20] , \edb_top_inst/la0/la_trig_mask[21] , 
        \edb_top_inst/la0/la_trig_mask[22] , \edb_top_inst/la0/la_trig_mask[23] , 
        \edb_top_inst/la0/la_trig_mask[24] , \edb_top_inst/la0/la_trig_mask[25] , 
        \edb_top_inst/la0/la_trig_mask[26] , \edb_top_inst/la0/la_trig_mask[27] , 
        \edb_top_inst/la0/la_trig_mask[28] , \edb_top_inst/la0/la_trig_mask[29] , 
        \edb_top_inst/la0/la_trig_mask[30] , \edb_top_inst/la0/la_trig_mask[31] , 
        \edb_top_inst/la0/la_trig_mask[32] , \edb_top_inst/la0/la_trig_mask[33] , 
        \edb_top_inst/la0/la_trig_mask[34] , \edb_top_inst/la0/la_trig_mask[35] , 
        \edb_top_inst/la0/la_trig_mask[36] , \edb_top_inst/la0/la_trig_mask[37] , 
        \edb_top_inst/la0/la_trig_mask[38] , \edb_top_inst/la0/la_trig_mask[39] , 
        \edb_top_inst/la0/la_trig_mask[40] , \edb_top_inst/la0/la_trig_mask[41] , 
        \edb_top_inst/la0/la_trig_mask[42] , \edb_top_inst/la0/la_trig_mask[43] , 
        \edb_top_inst/la0/la_trig_mask[44] , \edb_top_inst/la0/la_trig_mask[45] , 
        \edb_top_inst/la0/la_trig_mask[46] , \edb_top_inst/la0/la_trig_mask[47] , 
        \edb_top_inst/la0/la_trig_mask[48] , \edb_top_inst/la0/la_trig_mask[49] , 
        \edb_top_inst/la0/la_trig_mask[50] , \edb_top_inst/la0/la_trig_mask[51] , 
        \edb_top_inst/la0/la_trig_mask[52] , \edb_top_inst/la0/la_trig_mask[53] , 
        \edb_top_inst/la0/la_trig_mask[54] , \edb_top_inst/la0/la_trig_mask[55] , 
        \edb_top_inst/la0/la_trig_mask[56] , \edb_top_inst/la0/la_trig_mask[57] , 
        \edb_top_inst/la0/la_trig_mask[58] , \edb_top_inst/la0/la_trig_mask[59] , 
        \edb_top_inst/la0/la_trig_mask[60] , \edb_top_inst/la0/la_trig_mask[61] , 
        \edb_top_inst/la0/la_trig_mask[62] , \edb_top_inst/la0/la_trig_mask[63] , 
        \edb_top_inst/la0/la_num_trigger[1] , \edb_top_inst/la0/la_num_trigger[2] , 
        \edb_top_inst/la0/la_num_trigger[3] , \edb_top_inst/la0/la_num_trigger[4] , 
        \edb_top_inst/la0/la_num_trigger[5] , \edb_top_inst/la0/la_num_trigger[6] , 
        \edb_top_inst/la0/la_num_trigger[7] , \edb_top_inst/la0/la_num_trigger[8] , 
        \edb_top_inst/la0/la_num_trigger[9] , \edb_top_inst/la0/la_num_trigger[10] , 
        \edb_top_inst/la0/la_num_trigger[11] , \edb_top_inst/la0/la_num_trigger[12] , 
        \edb_top_inst/la0/la_num_trigger[13] , \edb_top_inst/la0/la_num_trigger[14] , 
        \edb_top_inst/la0/la_num_trigger[15] , \edb_top_inst/la0/la_num_trigger[16] , 
        \edb_top_inst/la0/la_window_depth[1] , \edb_top_inst/la0/la_window_depth[2] , 
        \edb_top_inst/la0/la_window_depth[3] , \edb_top_inst/la0/la_window_depth[4] , 
        \edb_top_inst/la0/address_counter[1] , \edb_top_inst/la0/address_counter[2] , 
        \edb_top_inst/la0/address_counter[3] , \edb_top_inst/la0/address_counter[4] , 
        \edb_top_inst/la0/address_counter[5] , \edb_top_inst/la0/address_counter[6] , 
        \edb_top_inst/la0/address_counter[7] , \edb_top_inst/la0/address_counter[8] , 
        \edb_top_inst/la0/address_counter[9] , \edb_top_inst/la0/address_counter[10] , 
        \edb_top_inst/la0/address_counter[11] , \edb_top_inst/la0/address_counter[12] , 
        \edb_top_inst/la0/address_counter[13] , \edb_top_inst/la0/address_counter[14] , 
        \edb_top_inst/la0/address_counter[15] , \edb_top_inst/la0/address_counter[16] , 
        \edb_top_inst/la0/address_counter[17] , \edb_top_inst/la0/address_counter[18] , 
        \edb_top_inst/la0/address_counter[19] , \edb_top_inst/la0/address_counter[20] , 
        \edb_top_inst/la0/address_counter[21] , \edb_top_inst/la0/address_counter[22] , 
        \edb_top_inst/la0/address_counter[23] , \edb_top_inst/la0/address_counter[24] , 
        \edb_top_inst/la0/address_counter[25] , \edb_top_inst/la0/opcode[1] , 
        \edb_top_inst/la0/opcode[2] , \edb_top_inst/la0/opcode[3] , \edb_top_inst/la0/bit_count[1] , 
        \edb_top_inst/la0/bit_count[2] , \edb_top_inst/la0/bit_count[3] , 
        \edb_top_inst/la0/bit_count[4] , \edb_top_inst/la0/bit_count[5] , 
        \edb_top_inst/la0/word_count[1] , \edb_top_inst/la0/word_count[2] , 
        \edb_top_inst/la0/word_count[3] , \edb_top_inst/la0/word_count[4] , 
        \edb_top_inst/la0/word_count[5] , \edb_top_inst/la0/word_count[6] , 
        \edb_top_inst/la0/word_count[7] , \edb_top_inst/la0/word_count[8] , 
        \edb_top_inst/la0/word_count[9] , \edb_top_inst/la0/word_count[10] , 
        \edb_top_inst/la0/word_count[11] , \edb_top_inst/la0/word_count[12] , 
        \edb_top_inst/la0/word_count[13] , \edb_top_inst/la0/word_count[14] , 
        \edb_top_inst/la0/word_count[15] , \edb_top_inst/la0/data_out_shift_reg[1] , 
        \edb_top_inst/la0/data_out_shift_reg[2] , \edb_top_inst/la0/data_out_shift_reg[3] , 
        \edb_top_inst/la0/data_out_shift_reg[4] , \edb_top_inst/la0/data_out_shift_reg[5] , 
        \edb_top_inst/la0/data_out_shift_reg[6] , \edb_top_inst/la0/data_out_shift_reg[7] , 
        \edb_top_inst/la0/data_out_shift_reg[8] , \edb_top_inst/la0/data_out_shift_reg[9] , 
        \edb_top_inst/la0/data_out_shift_reg[10] , \edb_top_inst/la0/data_out_shift_reg[11] , 
        \edb_top_inst/la0/data_out_shift_reg[12] , \edb_top_inst/la0/data_out_shift_reg[13] , 
        \edb_top_inst/la0/data_out_shift_reg[14] , \edb_top_inst/la0/data_out_shift_reg[15] , 
        \edb_top_inst/la0/data_out_shift_reg[16] , \edb_top_inst/la0/data_out_shift_reg[17] , 
        \edb_top_inst/la0/data_out_shift_reg[18] , \edb_top_inst/la0/data_out_shift_reg[19] , 
        \edb_top_inst/la0/data_out_shift_reg[20] , \edb_top_inst/la0/data_out_shift_reg[21] , 
        \edb_top_inst/la0/data_out_shift_reg[22] , \edb_top_inst/la0/data_out_shift_reg[23] , 
        \edb_top_inst/la0/data_out_shift_reg[24] , \edb_top_inst/la0/data_out_shift_reg[25] , 
        \edb_top_inst/la0/data_out_shift_reg[26] , \edb_top_inst/la0/data_out_shift_reg[27] , 
        \edb_top_inst/la0/data_out_shift_reg[28] , \edb_top_inst/la0/data_out_shift_reg[29] , 
        \edb_top_inst/la0/data_out_shift_reg[30] , \edb_top_inst/la0/data_out_shift_reg[31] , 
        \edb_top_inst/la0/data_out_shift_reg[32] , \edb_top_inst/la0/data_out_shift_reg[33] , 
        \edb_top_inst/la0/data_out_shift_reg[34] , \edb_top_inst/la0/data_out_shift_reg[35] , 
        \edb_top_inst/la0/data_out_shift_reg[36] , \edb_top_inst/la0/data_out_shift_reg[37] , 
        \edb_top_inst/la0/data_out_shift_reg[38] , \edb_top_inst/la0/data_out_shift_reg[39] , 
        \edb_top_inst/la0/data_out_shift_reg[40] , \edb_top_inst/la0/data_out_shift_reg[41] , 
        \edb_top_inst/la0/data_out_shift_reg[42] , \edb_top_inst/la0/data_out_shift_reg[43] , 
        \edb_top_inst/la0/data_out_shift_reg[44] , \edb_top_inst/la0/data_out_shift_reg[45] , 
        \edb_top_inst/la0/data_out_shift_reg[46] , \edb_top_inst/la0/data_out_shift_reg[47] , 
        \edb_top_inst/la0/data_out_shift_reg[48] , \edb_top_inst/la0/data_out_shift_reg[49] , 
        \edb_top_inst/la0/data_out_shift_reg[50] , \edb_top_inst/la0/data_out_shift_reg[51] , 
        \edb_top_inst/la0/data_out_shift_reg[52] , \edb_top_inst/la0/data_out_shift_reg[53] , 
        \edb_top_inst/la0/data_out_shift_reg[54] , \edb_top_inst/la0/data_out_shift_reg[55] , 
        \edb_top_inst/la0/data_out_shift_reg[56] , \edb_top_inst/la0/data_out_shift_reg[57] , 
        \edb_top_inst/la0/data_out_shift_reg[58] , \edb_top_inst/la0/data_out_shift_reg[59] , 
        \edb_top_inst/la0/data_out_shift_reg[60] , \edb_top_inst/la0/data_out_shift_reg[61] , 
        \edb_top_inst/la0/data_out_shift_reg[62] , \edb_top_inst/la0/data_out_shift_reg[63] , 
        \edb_top_inst/la0/module_state[1] , \edb_top_inst/la0/module_state[2] , 
        \edb_top_inst/la0/module_state[3] , \edb_top_inst/la0/crc_data_out[0] , 
        \edb_top_inst/la0/crc_data_out[1] , \edb_top_inst/la0/crc_data_out[2] , 
        \edb_top_inst/la0/crc_data_out[3] , \edb_top_inst/la0/crc_data_out[4] , 
        \edb_top_inst/la0/crc_data_out[5] , \edb_top_inst/la0/crc_data_out[6] , 
        \edb_top_inst/la0/crc_data_out[7] , \edb_top_inst/la0/crc_data_out[8] , 
        \edb_top_inst/la0/crc_data_out[9] , \edb_top_inst/la0/crc_data_out[10] , 
        \edb_top_inst/la0/crc_data_out[11] , \edb_top_inst/la0/crc_data_out[12] , 
        \edb_top_inst/la0/crc_data_out[13] , \edb_top_inst/la0/crc_data_out[14] , 
        \edb_top_inst/la0/crc_data_out[15] , \edb_top_inst/la0/crc_data_out[16] , 
        \edb_top_inst/la0/crc_data_out[17] , \edb_top_inst/la0/crc_data_out[18] , 
        \edb_top_inst/la0/crc_data_out[19] , \edb_top_inst/la0/crc_data_out[20] , 
        \edb_top_inst/la0/crc_data_out[21] , \edb_top_inst/la0/crc_data_out[22] , 
        \edb_top_inst/la0/crc_data_out[23] , \edb_top_inst/la0/crc_data_out[24] , 
        \edb_top_inst/la0/crc_data_out[25] , \edb_top_inst/la0/crc_data_out[26] , 
        \edb_top_inst/la0/crc_data_out[27] , \edb_top_inst/la0/crc_data_out[28] , 
        \edb_top_inst/la0/crc_data_out[29] , \edb_top_inst/la0/crc_data_out[30] , 
        \edb_top_inst/la0/crc_data_out[31] , \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.cap_probe_cout , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.cap_probe_cout , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9] , \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11] , \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13] , \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14] , 
        \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15] , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.cap_probe_cout , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[8] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[9] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[10] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[11] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[12] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[13] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[14] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[15] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] , \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.cap_probe_cout , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7] , 
        \edb_top_inst/la0/genblk2.la_capture_mask[1] , \edb_top_inst/la0/genblk2.la_capture_mask[2] , 
        \edb_top_inst/la0/genblk2.la_capture_mask[3] , \edb_top_inst/la0/genblk2.la_capture_mask[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.cap_probe_cout , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] , 
        \edb_top_inst/la0/tu_trigger , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26] , \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27] , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28] , \edb_top_inst/la0/capture_enable , 
        \edb_top_inst/la0/cap_fifo_din_cu[2] , \edb_top_inst/la0/cap_fifo_din_cu[3] , 
        \edb_top_inst/la0/cap_fifo_din_cu[4] , \edb_top_inst/la0/cap_fifo_din_cu[5] , 
        \edb_top_inst/la0/cap_fifo_din_cu[6] , \edb_top_inst/la0/cap_fifo_din_cu[7] , 
        \edb_top_inst/la0/cap_fifo_din_cu[8] , \edb_top_inst/la0/cap_fifo_din_cu[9] , 
        \edb_top_inst/la0/cap_fifo_din_cu[10] , \edb_top_inst/la0/cap_fifo_din_cu[11] , 
        \edb_top_inst/la0/cap_fifo_din_cu[12] , \edb_top_inst/la0/cap_fifo_din_cu[13] , 
        \edb_top_inst/la0/cap_fifo_din_cu[14] , \edb_top_inst/la0/cap_fifo_din_cu[15] , 
        \edb_top_inst/la0/cap_fifo_din_cu[16] , \edb_top_inst/la0/cap_fifo_din_cu[17] , 
        \edb_top_inst/la0/cap_fifo_din_cu[18] , \edb_top_inst/la0/cap_fifo_din_cu[19] , 
        \edb_top_inst/la0/cap_fifo_din_cu[20] , \edb_top_inst/la0/cap_fifo_din_cu[21] , 
        \edb_top_inst/la0/cap_fifo_din_cu[22] , \edb_top_inst/la0/cap_fifo_din_cu[23] , 
        \edb_top_inst/la0/cap_fifo_din_cu[24] , \edb_top_inst/la0/cap_fifo_din_cu[25] , 
        \edb_top_inst/la0/cap_fifo_din_cu[26] , \edb_top_inst/la0/cap_fifo_din_cu[27] , 
        \edb_top_inst/la0/cap_fifo_din_cu[28] , \edb_top_inst/la0/cap_fifo_din_tu[1] , 
        \edb_top_inst/la0/cap_fifo_din_tu[2] , \edb_top_inst/la0/cap_fifo_din_tu[3] , 
        \edb_top_inst/la0/cap_fifo_din_tu[4] , \edb_top_inst/la0/cap_fifo_din_tu[5] , 
        \edb_top_inst/la0/cap_fifo_din_tu[6] , \edb_top_inst/la0/cap_fifo_din_tu[7] , 
        \edb_top_inst/la0/cap_fifo_din_tu[8] , \edb_top_inst/la0/cap_fifo_din_tu[9] , 
        \edb_top_inst/la0/cap_fifo_din_tu[10] , \edb_top_inst/la0/cap_fifo_din_tu[11] , 
        \edb_top_inst/la0/cap_fifo_din_tu[12] , \edb_top_inst/la0/cap_fifo_din_tu[13] , 
        \edb_top_inst/la0/cap_fifo_din_tu[14] , \edb_top_inst/la0/cap_fifo_din_tu[15] , 
        \edb_top_inst/la0/cap_fifo_din_tu[16] , \edb_top_inst/la0/cap_fifo_din_tu[17] , 
        \edb_top_inst/la0/cap_fifo_din_tu[18] , \edb_top_inst/la0/cap_fifo_din_tu[19] , 
        \edb_top_inst/la0/cap_fifo_din_tu[20] , \edb_top_inst/la0/cap_fifo_din_tu[21] , 
        \edb_top_inst/la0/cap_fifo_din_tu[22] , \edb_top_inst/la0/cap_fifo_din_tu[23] , 
        \edb_top_inst/la0/cap_fifo_din_tu[24] , \edb_top_inst/la0/cap_fifo_din_tu[25] , 
        \edb_top_inst/la0/cap_fifo_din_tu[26] , \edb_top_inst/la0/cap_fifo_din_tu[27] , 
        \edb_top_inst/la0/cap_fifo_din_tu[28] , \edb_top_inst/la0/la_biu_inst/curr_state[0] , 
        \edb_top_inst/la0/la_biu_inst/run_trig_p2 , \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 , 
        \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 , \edb_top_inst/la0/la_biu_inst/str_sync , 
        \edb_top_inst/la0/la_biu_inst/str_sync_wbff1 , \edb_top_inst/la0/la_biu_inst/str_sync_wbff2 , 
        \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q , \edb_top_inst/la0/la_biu_inst/rdy_sync , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 , \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 , 
        \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q , \edb_top_inst/la0/data_from_biu[0] , 
        \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] , \edb_top_inst/la0/la_biu_inst/curr_state[3] , 
        \edb_top_inst/la0/la_biu_inst/curr_state[2] , \edb_top_inst/la0/la_biu_inst/curr_state[1] , 
        \edb_top_inst/la0/biu_ready , \edb_top_inst/la0/la_biu_inst/addr_reg[15] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[16] , \edb_top_inst/la0/la_biu_inst/addr_reg[17] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[18] , \edb_top_inst/la0/la_biu_inst/addr_reg[19] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[20] , \edb_top_inst/la0/la_biu_inst/addr_reg[21] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[22] , \edb_top_inst/la0/la_biu_inst/addr_reg[23] , 
        \edb_top_inst/la0/la_biu_inst/addr_reg[24] , \edb_top_inst/la0/la_biu_inst/addr_reg[25] , 
        \edb_top_inst/la0/data_from_biu[1] , \edb_top_inst/la0/data_from_biu[2] , 
        \edb_top_inst/la0/data_from_biu[3] , \edb_top_inst/la0/data_from_biu[4] , 
        \edb_top_inst/la0/data_from_biu[5] , \edb_top_inst/la0/data_from_biu[6] , 
        \edb_top_inst/la0/data_from_biu[7] , \edb_top_inst/la0/data_from_biu[8] , 
        \edb_top_inst/la0/data_from_biu[9] , \edb_top_inst/la0/data_from_biu[10] , 
        \edb_top_inst/la0/data_from_biu[11] , \edb_top_inst/la0/data_from_biu[12] , 
        \edb_top_inst/la0/data_from_biu[13] , \edb_top_inst/la0/data_from_biu[14] , 
        \edb_top_inst/la0/data_from_biu[15] , \edb_top_inst/la0/data_from_biu[16] , 
        \edb_top_inst/la0/data_from_biu[17] , \edb_top_inst/la0/data_from_biu[18] , 
        \edb_top_inst/la0/data_from_biu[19] , \edb_top_inst/la0/data_from_biu[20] , 
        \edb_top_inst/la0/data_from_biu[21] , \edb_top_inst/la0/data_from_biu[22] , 
        \edb_top_inst/la0/data_from_biu[23] , \edb_top_inst/la0/data_from_biu[24] , 
        \edb_top_inst/la0/data_from_biu[25] , \edb_top_inst/la0/data_from_biu[26] , 
        \edb_top_inst/la0/data_from_biu[27] , \edb_top_inst/la0/data_from_biu[28] , 
        \edb_top_inst/la0/data_from_biu[29] , \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] , 
        \edb_top_inst/la0/la_sample_cnt[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[0] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] , \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] , 
        \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] , 
        \edb_top_inst/la0/la_sample_cnt[1] , \edb_top_inst/la0/la_sample_cnt[2] , 
        \edb_top_inst/la0/la_sample_cnt[3] , \edb_top_inst/la0/la_sample_cnt[4] , 
        \edb_top_inst/la0/la_sample_cnt[5] , \edb_top_inst/la0/la_sample_cnt[6] , 
        \edb_top_inst/la0/la_sample_cnt[7] , \edb_top_inst/la0/la_sample_cnt[8] , 
        \edb_top_inst/la0/la_sample_cnt[9] , \edb_top_inst/la0/la_sample_cnt[10] , 
        \edb_top_inst/la0/la_sample_cnt[11] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[1] , \edb_top_inst/la0/la_biu_inst/fifo_counter[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[3] , \edb_top_inst/la0/la_biu_inst/fifo_counter[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[5] , \edb_top_inst/la0/la_biu_inst/fifo_counter[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[7] , \edb_top_inst/la0/la_biu_inst/fifo_counter[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_counter[9] , \edb_top_inst/la0/la_biu_inst/fifo_counter[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[11] , \edb_top_inst/la0/internal_register_select[1] , 
        \edb_top_inst/la0/internal_register_select[2] , \edb_top_inst/la0/internal_register_select[3] , 
        \edb_top_inst/la0/internal_register_select[4] , \edb_top_inst/la0/internal_register_select[5] , 
        \edb_top_inst/la0/internal_register_select[6] , \edb_top_inst/la0/internal_register_select[7] , 
        \edb_top_inst/la0/internal_register_select[8] , \edb_top_inst/la0/internal_register_select[9] , 
        \edb_top_inst/la0/internal_register_select[10] , \edb_top_inst/la0/internal_register_select[11] , 
        \edb_top_inst/la0/internal_register_select[12] , \edb_top_inst/la0/la_trig_pos[1] , 
        \edb_top_inst/la0/la_trig_pos[2] , \edb_top_inst/la0/la_trig_pos[3] , 
        \edb_top_inst/la0/la_trig_pos[4] , \edb_top_inst/la0/la_trig_pos[5] , 
        \edb_top_inst/la0/la_trig_pos[6] , \edb_top_inst/la0/la_trig_pos[7] , 
        \edb_top_inst/la0/la_trig_pos[8] , \edb_top_inst/la0/la_trig_pos[9] , 
        \edb_top_inst/la0/la_trig_pos[10] , \edb_top_inst/la0/la_trig_pos[11] , 
        \edb_top_inst/la0/la_trig_pos[12] , \edb_top_inst/la0/la_trig_pos[13] , 
        \edb_top_inst/la0/la_trig_pos[14] , \edb_top_inst/la0/la_trig_pos[15] , 
        \edb_top_inst/la0/la_trig_pos[16] , \edb_top_inst/debug_hub_inst/module_id_reg[0] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[1] , \edb_top_inst/debug_hub_inst/module_id_reg[2] , 
        \edb_top_inst/debug_hub_inst/module_id_reg[3] , \edb_top_inst/n54 , 
        \edb_top_inst/n56 , \edb_top_inst/n342 , \edb_top_inst/n775 , 
        \edb_top_inst/n777 , \edb_top_inst/n779 , \edb_top_inst/n781 , 
        \edb_top_inst/n2271 , \edb_top_inst/n2272 , \edb_top_inst/n2273 , 
        \edb_top_inst/n2274 , \edb_top_inst/n2275 , \edb_top_inst/n2276 , 
        \edb_top_inst/n2277 , \edb_top_inst/n2278 , \edb_top_inst/n2279 , 
        \edb_top_inst/n2280 , \edb_top_inst/n2281 , \edb_top_inst/n2282 , 
        \edb_top_inst/n2283 , \edb_top_inst/n2284 , \edb_top_inst/n2285 , 
        \edb_top_inst/n2286 , \edb_top_inst/n2287 , \edb_top_inst/n2288 , 
        \edb_top_inst/n2289 , \edb_top_inst/n2290 , \edb_top_inst/n2291 , 
        \edb_top_inst/n2292 , \edb_top_inst/n2293 , \edb_top_inst/n2294 , 
        \edb_top_inst/n2295 , \edb_top_inst/n2296 , \edb_top_inst/n2297 , 
        \edb_top_inst/n2298 , \edb_top_inst/n2299 , \edb_top_inst/n2247 , 
        \edb_top_inst/n2244 , \edb_top_inst/n2300 , \edb_top_inst/n2301 , 
        \edb_top_inst/n2302 , \edb_top_inst/n1285 , \edb_top_inst/n2303 , 
        \edb_top_inst/n2304 , \edb_top_inst/n2305 , \edb_top_inst/n2306 , 
        \edb_top_inst/n2307 , \edb_top_inst/n2308 , \edb_top_inst/n2309 , 
        \edb_top_inst/n2310 , \edb_top_inst/n2311 , \edb_top_inst/n2312 , 
        \edb_top_inst/n2313 , \edb_top_inst/n2314 , \edb_top_inst/n2315 , 
        \edb_top_inst/n2316 , \edb_top_inst/n2317 , \edb_top_inst/n2318 , 
        \edb_top_inst/n2319 , \edb_top_inst/n2320 , \edb_top_inst/n2321 , 
        \edb_top_inst/n2322 , \edb_top_inst/n2323 , \edb_top_inst/n2324 , 
        \edb_top_inst/n2325 , \edb_top_inst/n2326 , \edb_top_inst/n2327 , 
        \edb_top_inst/n2328 , \edb_top_inst/n2329 , \edb_top_inst/n2330 , 
        \edb_top_inst/n2331 , \edb_top_inst/n2332 , \edb_top_inst/n2333 , 
        \edb_top_inst/n2334 , \edb_top_inst/n2335 , \edb_top_inst/n2336 , 
        \edb_top_inst/n2337 , \edb_top_inst/n2338 , \edb_top_inst/n2339 , 
        \edb_top_inst/n2340 , \edb_top_inst/n2341 , \edb_top_inst/n2342 , 
        \edb_top_inst/n2343 , \edb_top_inst/n2344 , \edb_top_inst/n2345 , 
        \edb_top_inst/n2346 , \edb_top_inst/n2347 , \edb_top_inst/n2348 , 
        \edb_top_inst/n2349 , \edb_top_inst/n2350 , \edb_top_inst/n2351 , 
        \edb_top_inst/n2352 , \edb_top_inst/n2353 , \edb_top_inst/n2354 , 
        \edb_top_inst/n2355 , \edb_top_inst/n2356 , \edb_top_inst/n2357 , 
        \edb_top_inst/n2358 , \edb_top_inst/n2359 , \edb_top_inst/n2360 , 
        \edb_top_inst/n2361 , \edb_top_inst/n2362 , \edb_top_inst/n2363 , 
        \edb_top_inst/n2364 , \edb_top_inst/n2365 , \edb_top_inst/n2366 , 
        \edb_top_inst/n2367 , \edb_top_inst/n2368 , \edb_top_inst/n2369 , 
        \edb_top_inst/n2370 , \edb_top_inst/n2371 , \edb_top_inst/n2372 , 
        \edb_top_inst/n2373 , \edb_top_inst/n2374 , \edb_top_inst/n2375 , 
        \edb_top_inst/n2376 , \edb_top_inst/n2377 , \edb_top_inst/n2378 , 
        \edb_top_inst/n2379 , \edb_top_inst/n2380 , \edb_top_inst/n2381 , 
        \edb_top_inst/n2382 , \edb_top_inst/n2383 , \edb_top_inst/n2384 , 
        \edb_top_inst/n2385 , \edb_top_inst/n2386 , \edb_top_inst/n2387 , 
        \edb_top_inst/n2388 , \edb_top_inst/n2389 , \edb_top_inst/n2390 , 
        \edb_top_inst/n2391 , \edb_top_inst/n2392 , \edb_top_inst/n2393 , 
        \edb_top_inst/n2394 , \edb_top_inst/n2401 , \edb_top_inst/n2402 , 
        \edb_top_inst/n2403 , \edb_top_inst/n2404 , \edb_top_inst/n2405 , 
        \edb_top_inst/n2406 , \edb_top_inst/n2407 , \edb_top_inst/n2408 , 
        \edb_top_inst/n2409 , \edb_top_inst/n2410 , \edb_top_inst/n2411 , 
        \edb_top_inst/n2412 , \edb_top_inst/n2413 , \edb_top_inst/n2414 , 
        \edb_top_inst/n2415 , \edb_top_inst/n2416 , \edb_top_inst/n2417 , 
        \edb_top_inst/n2418 , \edb_top_inst/n2419 , \edb_top_inst/n2420 , 
        \edb_top_inst/n2421 , \edb_top_inst/n2422 , \edb_top_inst/n2424 , 
        \edb_top_inst/n2425 , \edb_top_inst/n2426 , \edb_top_inst/n2427 , 
        \edb_top_inst/n2428 , \edb_top_inst/n2429 , \edb_top_inst/n2430 , 
        \edb_top_inst/n2431 , \edb_top_inst/n2432 , \edb_top_inst/n2433 , 
        \edb_top_inst/n2434 , \edb_top_inst/n2435 , \edb_top_inst/n2436 , 
        \edb_top_inst/n2437 , \edb_top_inst/n2438 , \edb_top_inst/n2439 , 
        \edb_top_inst/n2440 , \edb_top_inst/n2441 , \edb_top_inst/n2442 , 
        \edb_top_inst/n2443 , \edb_top_inst/n2444 , \edb_top_inst/n2445 , 
        \edb_top_inst/n2446 , \edb_top_inst/n2447 , \edb_top_inst/n2448 , 
        \edb_top_inst/n2449 , \edb_top_inst/n2450 , \edb_top_inst/n2451 , 
        \edb_top_inst/n2452 , \edb_top_inst/n2453 , \edb_top_inst/n2454 , 
        \edb_top_inst/n2455 , \edb_top_inst/n2456 , \edb_top_inst/n2457 , 
        \edb_top_inst/n2458 , \edb_top_inst/n2459 , \edb_top_inst/n2460 , 
        \edb_top_inst/n2461 , \edb_top_inst/n2462 , \edb_top_inst/n2463 , 
        \edb_top_inst/n2464 , \edb_top_inst/n2465 , \edb_top_inst/n2466 , 
        \edb_top_inst/n2467 , \edb_top_inst/n2468 , \edb_top_inst/n2469 , 
        \edb_top_inst/n2470 , \edb_top_inst/n2471 , \edb_top_inst/n2472 , 
        \edb_top_inst/n2473 , \edb_top_inst/n2474 , \edb_top_inst/n2475 , 
        \edb_top_inst/n2476 , \edb_top_inst/n2477 , \edb_top_inst/n2478 , 
        \edb_top_inst/n2479 , \edb_top_inst/n2480 , \edb_top_inst/n2481 , 
        \edb_top_inst/n2482 , \edb_top_inst/n2483 , \edb_top_inst/n2484 , 
        \edb_top_inst/n2485 , \edb_top_inst/n2486 , \edb_top_inst/n2487 , 
        \edb_top_inst/n2488 , \edb_top_inst/n2489 , \edb_top_inst/n2490 , 
        \edb_top_inst/n2491 , \edb_top_inst/n2492 , \edb_top_inst/n2493 , 
        \edb_top_inst/n2494 , \edb_top_inst/n2495 , \edb_top_inst/n2496 , 
        \edb_top_inst/n2497 , \edb_top_inst/n2498 , \edb_top_inst/n2499 , 
        \edb_top_inst/n2500 , \edb_top_inst/n2501 , \edb_top_inst/n2502 , 
        \edb_top_inst/n2503 , \edb_top_inst/n2504 , \edb_top_inst/n2505 , 
        \edb_top_inst/n2506 , \edb_top_inst/n2507 , \edb_top_inst/n2508 , 
        \edb_top_inst/n2509 , \edb_top_inst/n2510 , \edb_top_inst/n2511 , 
        \edb_top_inst/n2512 , \edb_top_inst/n2513 , \edb_top_inst/n2514 , 
        \edb_top_inst/n2515 , \edb_top_inst/n2516 , \edb_top_inst/n2517 , 
        \edb_top_inst/n2518 , \edb_top_inst/n2519 , \edb_top_inst/n2520 , 
        \edb_top_inst/n2521 , \edb_top_inst/n2522 , \edb_top_inst/n2523 , 
        \edb_top_inst/n2524 , \edb_top_inst/n2525 , \edb_top_inst/n2526 , 
        \edb_top_inst/n2527 , \edb_top_inst/n2528 , \edb_top_inst/n2529 , 
        \edb_top_inst/n2530 , \edb_top_inst/n2531 , \edb_top_inst/n2532 , 
        \edb_top_inst/n2533 , \edb_top_inst/n2534 , \edb_top_inst/n2535 , 
        \edb_top_inst/n2536 , \edb_top_inst/n2537 , \edb_top_inst/n2538 , 
        \edb_top_inst/n2539 , \edb_top_inst/n2540 , \edb_top_inst/n2541 , 
        \edb_top_inst/n2542 , \edb_top_inst/n2543 , \edb_top_inst/n2544 , 
        \edb_top_inst/n2545 , \edb_top_inst/n2546 , \edb_top_inst/n2547 , 
        \edb_top_inst/n2548 , \edb_top_inst/n2549 , \edb_top_inst/n2550 , 
        \edb_top_inst/n2551 , \edb_top_inst/n2552 , \edb_top_inst/n2553 , 
        \edb_top_inst/n2554 , \edb_top_inst/n2555 , \edb_top_inst/n2556 , 
        \edb_top_inst/n2557 , \edb_top_inst/n2558 , \edb_top_inst/n2559 , 
        \edb_top_inst/n2560 , \edb_top_inst/n2561 , \edb_top_inst/n2562 , 
        \edb_top_inst/n2563 , \edb_top_inst/n2564 , \edb_top_inst/n2565 , 
        \edb_top_inst/n2566 , \edb_top_inst/n2567 , \edb_top_inst/n2568 , 
        \edb_top_inst/n2569 , \edb_top_inst/n2570 , \edb_top_inst/n2571 , 
        \edb_top_inst/n2572 , \edb_top_inst/n2573 , \edb_top_inst/n2574 , 
        \edb_top_inst/n2575 , \edb_top_inst/n2576 , \edb_top_inst/n2577 , 
        \edb_top_inst/n2578 , \edb_top_inst/n2579 , \edb_top_inst/n2580 , 
        \edb_top_inst/n2581 , \edb_top_inst/n2582 , \edb_top_inst/n2583 , 
        \edb_top_inst/n2584 , \edb_top_inst/n2585 , \edb_top_inst/n2586 , 
        \edb_top_inst/n2587 , \edb_top_inst/n2588 , \edb_top_inst/n2589 , 
        \edb_top_inst/n2590 , \edb_top_inst/n2591 , \edb_top_inst/n2592 , 
        \edb_top_inst/n2593 , \edb_top_inst/n2594 , \edb_top_inst/n2595 , 
        \edb_top_inst/n2596 , \edb_top_inst/n2597 , \edb_top_inst/n2598 , 
        \edb_top_inst/n2599 , \edb_top_inst/n2600 , \edb_top_inst/n2601 , 
        \edb_top_inst/n2602 , \edb_top_inst/n2603 , \edb_top_inst/n2604 , 
        \edb_top_inst/n2605 , \edb_top_inst/n2606 , \edb_top_inst/n2607 , 
        \edb_top_inst/n2608 , \edb_top_inst/n2609 , \edb_top_inst/n2610 , 
        \edb_top_inst/n2611 , \edb_top_inst/n2612 , \edb_top_inst/n2613 , 
        \edb_top_inst/n2614 , \edb_top_inst/n2615 , \edb_top_inst/n2616 , 
        \edb_top_inst/n2617 , \edb_top_inst/n2618 , \edb_top_inst/n2619 , 
        \edb_top_inst/n2620 , \edb_top_inst/n2621 , \edb_top_inst/n2622 , 
        \edb_top_inst/n2623 , \edb_top_inst/n2624 , \edb_top_inst/n2625 , 
        \edb_top_inst/n2626 , \edb_top_inst/n2627 , \edb_top_inst/n2628 , 
        \edb_top_inst/n2629 , \edb_top_inst/n2630 , \edb_top_inst/n2631 , 
        \edb_top_inst/n2632 , \edb_top_inst/n2633 , \edb_top_inst/n2634 , 
        \edb_top_inst/n2635 , \edb_top_inst/n2636 , \edb_top_inst/n2637 , 
        \edb_top_inst/n2638 , \edb_top_inst/n2639 , \edb_top_inst/n2640 , 
        \edb_top_inst/n2641 , \edb_top_inst/n2642 , \edb_top_inst/n2643 , 
        \edb_top_inst/n2644 , \edb_top_inst/n2645 , \edb_top_inst/n2646 , 
        \edb_top_inst/n2647 , \edb_top_inst/n2648 , \edb_top_inst/n2649 , 
        \edb_top_inst/n2650 , \edb_top_inst/n2651 , \edb_top_inst/n2652 , 
        \edb_top_inst/n2653 , \edb_top_inst/n2654 , \edb_top_inst/n2655 , 
        \edb_top_inst/n2656 , \edb_top_inst/n2657 , \edb_top_inst/n2658 , 
        \edb_top_inst/n2659 , \edb_top_inst/n2660 , \edb_top_inst/n2661 , 
        \edb_top_inst/n2662 , \edb_top_inst/n2663 , \edb_top_inst/n2664 , 
        \edb_top_inst/n2665 , \edb_top_inst/n2666 , \edb_top_inst/n2667 , 
        \edb_top_inst/n2668 , \edb_top_inst/n2669 , \edb_top_inst/n2670 , 
        \edb_top_inst/n2671 , \edb_top_inst/n2672 , \edb_top_inst/n2673 , 
        \edb_top_inst/n2674 , \edb_top_inst/n2675 , \edb_top_inst/n2676 , 
        \edb_top_inst/n2677 , \edb_top_inst/n2678 , \edb_top_inst/n2679 , 
        \edb_top_inst/n2680 , \edb_top_inst/n2681 , \edb_top_inst/n2682 , 
        \edb_top_inst/n2683 , \edb_top_inst/n2684 , \edb_top_inst/n2685 , 
        \edb_top_inst/n2686 , \edb_top_inst/n2687 , \edb_top_inst/n2688 , 
        \edb_top_inst/n2689 , \edb_top_inst/n2690 , \edb_top_inst/n2691 , 
        \edb_top_inst/n2692 , \edb_top_inst/n2693 , \edb_top_inst/n2694 , 
        \edb_top_inst/n2695 , \edb_top_inst/n2696 , \edb_top_inst/n2697 , 
        \edb_top_inst/n2698 , \edb_top_inst/n2699 , \edb_top_inst/n2700 , 
        \edb_top_inst/n2701 , \edb_top_inst/n2702 , \edb_top_inst/n2703 , 
        \edb_top_inst/n2704 , \edb_top_inst/n2705 , \edb_top_inst/n2706 , 
        \edb_top_inst/n2707 , \edb_top_inst/n2708 , \edb_top_inst/n2709 , 
        \edb_top_inst/n2710 , \edb_top_inst/n2711 , \edb_top_inst/n2712 , 
        \edb_top_inst/n2713 , \edb_top_inst/n2714 , \edb_top_inst/n2715 , 
        \edb_top_inst/n2716 , \edb_top_inst/n2717 , \edb_top_inst/n2718 , 
        \edb_top_inst/n2719 , \edb_top_inst/n2720 , \edb_top_inst/n2721 , 
        \edb_top_inst/n2722 , \edb_top_inst/n2723 , \edb_top_inst/n2724 , 
        \edb_top_inst/n2725 , \edb_top_inst/n2726 , \edb_top_inst/n2727 , 
        \edb_top_inst/n2728 , \edb_top_inst/n2729 , \edb_top_inst/n2730 , 
        \edb_top_inst/n2731 , \edb_top_inst/n2732 , \edb_top_inst/n2733 , 
        \edb_top_inst/n2734 , \edb_top_inst/n2735 , \edb_top_inst/n2736 , 
        \edb_top_inst/n2737 , \edb_top_inst/n2738 , \edb_top_inst/n2739 , 
        \edb_top_inst/n2740 , \edb_top_inst/n2741 , \edb_top_inst/n2742 , 
        \edb_top_inst/n2743 , \edb_top_inst/n2744 , \edb_top_inst/n2745 , 
        \edb_top_inst/n2746 , \edb_top_inst/n2747 , \edb_top_inst/n2748 , 
        \edb_top_inst/n2749 , \edb_top_inst/n2750 , \edb_top_inst/n2751 , 
        \edb_top_inst/n2752 , \edb_top_inst/n2753 , \edb_top_inst/n2754 , 
        \edb_top_inst/n2755 , \edb_top_inst/n2756 , \edb_top_inst/n2757 , 
        \edb_top_inst/n2758 , \edb_top_inst/n2759 , \edb_top_inst/n2760 , 
        \edb_top_inst/n2761 , \edb_top_inst/n2762 , \edb_top_inst/n2763 , 
        \edb_top_inst/n2764 , \edb_top_inst/n2765 , \edb_top_inst/n2766 , 
        \edb_top_inst/n2767 , \edb_top_inst/n2768 , \edb_top_inst/n2769 , 
        \edb_top_inst/n2770 , \edb_top_inst/n2771 , \edb_top_inst/n2772 , 
        \edb_top_inst/n2773 , \edb_top_inst/n2774 , \edb_top_inst/n2775 , 
        \edb_top_inst/n2776 , \edb_top_inst/n2777 , \edb_top_inst/n2778 , 
        \edb_top_inst/n2779 , \edb_top_inst/n2780 , \edb_top_inst/n2781 , 
        \edb_top_inst/n2782 , \edb_top_inst/n2783 , \edb_top_inst/n2784 , 
        \edb_top_inst/n2785 , \edb_top_inst/n2786 , \edb_top_inst/n2787 , 
        \edb_top_inst/n2788 , \edb_top_inst/n2789 , \edb_top_inst/n2790 , 
        \edb_top_inst/n2791 , \edb_top_inst/n2792 , \edb_top_inst/n2793 , 
        \edb_top_inst/n2794 , \edb_top_inst/n2795 , \edb_top_inst/n2796 , 
        \edb_top_inst/n2797 , \edb_top_inst/n2798 , \edb_top_inst/n2799 , 
        \edb_top_inst/n2800 , \edb_top_inst/n2801 , \edb_top_inst/n2802 , 
        \edb_top_inst/n2803 , \edb_top_inst/n2804 , \edb_top_inst/n2805 , 
        \edb_top_inst/n2806 , \edb_top_inst/n2807 , \edb_top_inst/n2808 , 
        \edb_top_inst/n2809 , \edb_top_inst/n2810 , \edb_top_inst/n2811 , 
        \edb_top_inst/n2812 , \edb_top_inst/n2813 , \edb_top_inst/n2814 , 
        \edb_top_inst/n2815 , \edb_top_inst/n2816 , \edb_top_inst/n2817 , 
        \edb_top_inst/n2818 , \edb_top_inst/n2819 , \edb_top_inst/n2820 , 
        \edb_top_inst/n2821 , \edb_top_inst/n2822 , \edb_top_inst/n2823 , 
        \edb_top_inst/n2824 , \edb_top_inst/n2825 , \edb_top_inst/n2826 , 
        \edb_top_inst/n2827 , \edb_top_inst/n2828 , \edb_top_inst/n2829 , 
        \edb_top_inst/n2830 , \edb_top_inst/n2831 , \edb_top_inst/n2832 , 
        \edb_top_inst/n2833 , \edb_top_inst/n2834 , \edb_top_inst/n2835 , 
        \edb_top_inst/n2836 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , \edb_top_inst/n2837 , 
        \edb_top_inst/n2838 , \edb_top_inst/n2839 , \edb_top_inst/n2840 , 
        \edb_top_inst/n2841 , \edb_top_inst/n2842 , \edb_top_inst/n2843 , 
        \edb_top_inst/n2844 , \edb_top_inst/n2845 , \edb_top_inst/n2846 , 
        \edb_top_inst/n2847 , \edb_top_inst/n2848 , \edb_top_inst/n2849 , 
        \edb_top_inst/n2850 , \edb_top_inst/n2851 , \edb_top_inst/n2852 , 
        \edb_top_inst/n2853 , \edb_top_inst/n2854 , \edb_top_inst/n2855 , 
        \edb_top_inst/n2856 , \edb_top_inst/n2857 , \edb_top_inst/n2858 , 
        \edb_top_inst/n2859 , \edb_top_inst/n2860 , \edb_top_inst/n2861 , 
        \edb_top_inst/n2862 , \edb_top_inst/n2863 , \edb_top_inst/n2864 , 
        \edb_top_inst/n2865 , \edb_top_inst/n2866 , \edb_top_inst/n2867 , 
        \edb_top_inst/n2868 , \edb_top_inst/n2869 , \edb_top_inst/n2870 , 
        \edb_top_inst/n2871 , \edb_top_inst/n2872 , \edb_top_inst/n2873 , 
        \edb_top_inst/n2874 , \edb_top_inst/n2875 , \edb_top_inst/n2876 , 
        \edb_top_inst/n2877 , \edb_top_inst/n2878 , \edb_top_inst/n2250 , 
        \received_data[0] , ceg_net98, \state[1] , ceg_net127, \state[0] , 
        ceg_net130, ceg_net133, ceg_net108, \equal_4/n3 , ceg_net120, 
        ceg_net138, \uart_rx/n375 , ceg_net78, \uart_rx/n407 , ceg_net153, 
        \uart_rx/n444 , \uart_rx/n382 , ceg_net146, \uart_rx/n372 , 
        \uart_rx/r_SM_Main[2] , \uart_rx/n316 , \uart_rx/n319 , \uart_rx/n322 , 
        \uart_rx/n325 , \uart_rx/n328 , \uart_rx/n331 , \uart_rx/n334 , 
        \uart_rx/n429 , \uart_rx/n431 , \uart_rx/n433 , \uart_rx/n435 , 
        \uart_rx/n437 , \uart_rx/n439 , \uart_rx/n441 , \uart_rx/n359 , 
        \uart_rx/n363 , \uart_rx/n309 , \uart_rx/n43 , \uart_rx/n385 , 
        \received_data[1] , \received_data[2] , \received_data[3] , \received_data[4] , 
        \received_data[5] , \received_data[6] , \received_data[7] , n57, 
        \equal_5/n3 , \uart_tx1/n119 , \uart_tx1/n110 , \uart_tx1/select_38/Select_0/n3 , 
        \data_to_transmitter[0] , \uart_tx1/n338 , \uart_tx1/n138 , \uart_tx1/n118 , 
        \uart_tx1/n117 , \uart_tx1/n116 , \uart_tx1/n115 , \uart_tx1/n114 , 
        \uart_tx1/n113 , \uart_tx1/n122 , \uart_tx1/n121 , \data_to_transmitter[1] , 
        \data_to_transmitter[2] , \data_to_transmitter[3] , \data_to_transmitter[4] , 
        \data_to_transmitter[5] , \data_to_transmitter[6] , \data_to_transmitter[7] , 
        \uart_tx1/n137 , \uart_tx2/n110 , \data_to_transmitter[8] , \data_to_transmitter[9] , 
        \data_to_transmitter[10] , \data_to_transmitter[11] , \data_to_transmitter[12] , 
        \data_to_transmitter[13] , \data_to_transmitter[14] , \data_to_transmitter[15] , 
        \edb_top_inst/edb_user_dr[50] , \edb_top_inst/edb_user_dr[51] , 
        \edb_top_inst/la0/n1334 , \edb_top_inst/ceg_net5 , \edb_top_inst/edb_user_dr[60] , 
        \edb_top_inst/la0/n1306 , \edb_top_inst/la0/n1335 , \edb_top_inst/la0/n1336 , 
        \edb_top_inst/edb_user_dr[62] , \edb_top_inst/edb_user_dr[0] , \edb_top_inst/la0/n1390 , 
        \edb_top_inst/edb_user_dr[42] , \edb_top_inst/la0/n1907 , \edb_top_inst/edb_user_dr[59] , 
        \edb_top_inst/la0/n1959 , \edb_top_inst/la0/data_to_addr_counter[0] , 
        \edb_top_inst/la0/addr_ct_en , \edb_top_inst/edb_user_dr[77] , \edb_top_inst/la0/op_reg_en , 
        \edb_top_inst/la0/n2183 , \edb_top_inst/ceg_net26 , \edb_top_inst/la0/data_to_word_counter[0] , 
        \edb_top_inst/la0/word_ct_en , \edb_top_inst/la0/n2460 , \edb_top_inst/ceg_net14 , 
        \edb_top_inst/la0/module_next_state[0] , \edb_top_inst/la0/n2774 , 
        \edb_top_inst/la0/n2789 , \edb_top_inst/la0/n2987 , \edb_top_inst/la0/n3185 , 
        \edb_top_inst/la0/n3200 , \edb_top_inst/la0/n3398 , \edb_top_inst/edb_user_dr[1] , 
        \edb_top_inst/la0/n3611 , \edb_top_inst/la0/n4022 , \edb_top_inst/la0/n4460 , 
        \edb_top_inst/la0/n4475 , \edb_top_inst/la0/n4673 , \edb_top_inst/la0/n4871 , 
        \edb_top_inst/la0/n4886 , \edb_top_inst/la0/n5084 , \edb_top_inst/la0/n5409 , 
        \edb_top_inst/la0/n5424 , \edb_top_inst/la0/n5622 , \edb_top_inst/la0/n5820 , 
        \edb_top_inst/la0/n5835 , \edb_top_inst/la0/n6033 , \edb_top_inst/la0/n6316 , 
        \edb_top_inst/la0/n6331 , \edb_top_inst/la0/n6529 , \edb_top_inst/la0/n6727 , 
        \edb_top_inst/la0/n6742 , \edb_top_inst/la0/n6940 , \edb_top_inst/la0/n7152 , 
        \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1] , \edb_top_inst/edb_user_dr[64] , 
        \edb_top_inst/la0/regsel_ld_en , \edb_top_inst/edb_user_dr[43] , 
        \edb_top_inst/edb_user_dr[61] , \edb_top_inst/edb_user_dr[63] , 
        \edb_top_inst/edb_user_dr[2] , \edb_top_inst/edb_user_dr[3] , \edb_top_inst/edb_user_dr[4] , 
        \edb_top_inst/edb_user_dr[5] , \edb_top_inst/edb_user_dr[6] , \edb_top_inst/edb_user_dr[7] , 
        \edb_top_inst/edb_user_dr[8] , \edb_top_inst/edb_user_dr[9] , \edb_top_inst/edb_user_dr[10] , 
        \edb_top_inst/edb_user_dr[11] , \edb_top_inst/edb_user_dr[12] , 
        \edb_top_inst/edb_user_dr[13] , \edb_top_inst/edb_user_dr[14] , 
        \edb_top_inst/edb_user_dr[15] , \edb_top_inst/edb_user_dr[16] , 
        \edb_top_inst/edb_user_dr[17] , \edb_top_inst/edb_user_dr[18] , 
        \edb_top_inst/edb_user_dr[19] , \edb_top_inst/edb_user_dr[20] , 
        \edb_top_inst/edb_user_dr[21] , \edb_top_inst/edb_user_dr[22] , 
        \edb_top_inst/edb_user_dr[23] , \edb_top_inst/edb_user_dr[24] , 
        \edb_top_inst/edb_user_dr[25] , \edb_top_inst/edb_user_dr[26] , 
        \edb_top_inst/edb_user_dr[27] , \edb_top_inst/edb_user_dr[28] , 
        \edb_top_inst/edb_user_dr[29] , \edb_top_inst/edb_user_dr[30] , 
        \edb_top_inst/edb_user_dr[31] , \edb_top_inst/edb_user_dr[32] , 
        \edb_top_inst/edb_user_dr[33] , \edb_top_inst/edb_user_dr[34] , 
        \edb_top_inst/edb_user_dr[35] , \edb_top_inst/edb_user_dr[36] , 
        \edb_top_inst/edb_user_dr[37] , \edb_top_inst/edb_user_dr[38] , 
        \edb_top_inst/edb_user_dr[39] , \edb_top_inst/edb_user_dr[40] , 
        \edb_top_inst/edb_user_dr[41] , \edb_top_inst/edb_user_dr[44] , 
        \edb_top_inst/edb_user_dr[45] , \edb_top_inst/edb_user_dr[46] , 
        \edb_top_inst/edb_user_dr[47] , \edb_top_inst/edb_user_dr[48] , 
        \edb_top_inst/edb_user_dr[49] , \edb_top_inst/edb_user_dr[52] , 
        \edb_top_inst/edb_user_dr[53] , \edb_top_inst/edb_user_dr[54] , 
        \edb_top_inst/edb_user_dr[55] , \edb_top_inst/edb_user_dr[56] , 
        \edb_top_inst/edb_user_dr[57] , \edb_top_inst/edb_user_dr[58] , 
        \edb_top_inst/la0/data_to_addr_counter[1] , \edb_top_inst/la0/data_to_addr_counter[2] , 
        \edb_top_inst/la0/data_to_addr_counter[3] , \edb_top_inst/la0/data_to_addr_counter[4] , 
        \edb_top_inst/la0/data_to_addr_counter[5] , \edb_top_inst/la0/data_to_addr_counter[6] , 
        \edb_top_inst/la0/data_to_addr_counter[7] , \edb_top_inst/la0/data_to_addr_counter[8] , 
        \edb_top_inst/la0/data_to_addr_counter[9] , \edb_top_inst/la0/data_to_addr_counter[10] , 
        \edb_top_inst/la0/data_to_addr_counter[11] , \edb_top_inst/la0/data_to_addr_counter[12] , 
        \edb_top_inst/la0/data_to_addr_counter[13] , \edb_top_inst/la0/data_to_addr_counter[14] , 
        \edb_top_inst/la0/data_to_addr_counter[15] , \edb_top_inst/la0/data_to_addr_counter[16] , 
        \edb_top_inst/la0/data_to_addr_counter[17] , \edb_top_inst/la0/data_to_addr_counter[18] , 
        \edb_top_inst/la0/data_to_addr_counter[19] , \edb_top_inst/la0/data_to_addr_counter[20] , 
        \edb_top_inst/la0/data_to_addr_counter[21] , \edb_top_inst/la0/data_to_addr_counter[22] , 
        \edb_top_inst/la0/data_to_addr_counter[23] , \edb_top_inst/la0/data_to_addr_counter[24] , 
        \edb_top_inst/la0/data_to_addr_counter[25] , \edb_top_inst/edb_user_dr[78] , 
        \edb_top_inst/edb_user_dr[79] , \edb_top_inst/edb_user_dr[80] , 
        \edb_top_inst/la0/n2182 , \edb_top_inst/la0/n2181 , \edb_top_inst/la0/n2180 , 
        \edb_top_inst/la0/n2179 , \edb_top_inst/la0/n2178 , \edb_top_inst/la0/data_to_word_counter[1] , 
        \edb_top_inst/la0/data_to_word_counter[2] , \edb_top_inst/la0/data_to_word_counter[3] , 
        \edb_top_inst/la0/data_to_word_counter[4] , \edb_top_inst/la0/data_to_word_counter[5] , 
        \edb_top_inst/la0/data_to_word_counter[6] , \edb_top_inst/la0/data_to_word_counter[7] , 
        \edb_top_inst/la0/data_to_word_counter[8] , \edb_top_inst/la0/data_to_word_counter[9] , 
        \edb_top_inst/la0/data_to_word_counter[10] , \edb_top_inst/la0/data_to_word_counter[11] , 
        \edb_top_inst/la0/data_to_word_counter[12] , \edb_top_inst/la0/data_to_word_counter[13] , 
        \edb_top_inst/la0/data_to_word_counter[14] , \edb_top_inst/la0/data_to_word_counter[15] , 
        \edb_top_inst/la0/n2459 , \edb_top_inst/la0/n2458 , \edb_top_inst/la0/n2457 , 
        \edb_top_inst/la0/n2456 , \edb_top_inst/la0/n2455 , \edb_top_inst/la0/n2454 , 
        \edb_top_inst/la0/n2453 , \edb_top_inst/la0/n2452 , \edb_top_inst/la0/n2451 , 
        \edb_top_inst/la0/n2450 , \edb_top_inst/la0/n2449 , \edb_top_inst/la0/n2448 , 
        \edb_top_inst/la0/n2447 , \edb_top_inst/la0/n2446 , \edb_top_inst/la0/n2445 , 
        \edb_top_inst/la0/n2444 , \edb_top_inst/la0/n2443 , \edb_top_inst/la0/n2442 , 
        \edb_top_inst/la0/n2441 , \edb_top_inst/la0/n2440 , \edb_top_inst/la0/n2439 , 
        \edb_top_inst/la0/n2438 , \edb_top_inst/la0/n2437 , \edb_top_inst/la0/n2436 , 
        \edb_top_inst/la0/n2435 , \edb_top_inst/la0/n2434 , \edb_top_inst/la0/n2433 , 
        \edb_top_inst/la0/n2432 , \edb_top_inst/la0/n2431 , \edb_top_inst/la0/n2430 , 
        \edb_top_inst/la0/n2429 , \edb_top_inst/la0/n2428 , \edb_top_inst/la0/n2427 , 
        \edb_top_inst/la0/n2426 , \edb_top_inst/la0/n2425 , \edb_top_inst/la0/n2424 , 
        \edb_top_inst/la0/n2423 , \edb_top_inst/la0/n2422 , \edb_top_inst/la0/n2421 , 
        \edb_top_inst/la0/n2420 , \edb_top_inst/la0/n2419 , \edb_top_inst/la0/n2418 , 
        \edb_top_inst/la0/n2417 , \edb_top_inst/la0/n2416 , \edb_top_inst/la0/n2415 , 
        \edb_top_inst/la0/n2414 , \edb_top_inst/la0/n2413 , \edb_top_inst/la0/n2412 , 
        \edb_top_inst/la0/n2411 , \edb_top_inst/la0/n2410 , \edb_top_inst/la0/n2409 , 
        \edb_top_inst/la0/n2408 , \edb_top_inst/la0/n2407 , \edb_top_inst/la0/n2406 , 
        \edb_top_inst/la0/n2405 , \edb_top_inst/la0/n2404 , \edb_top_inst/la0/n2403 , 
        \edb_top_inst/la0/n2402 , \edb_top_inst/la0/n2401 , \edb_top_inst/la0/n2400 , 
        \edb_top_inst/la0/n2399 , \edb_top_inst/la0/n2398 , \edb_top_inst/la0/n2397 , 
        \edb_top_inst/la0/module_next_state[1] , \edb_top_inst/la0/module_next_state[2] , 
        \edb_top_inst/la0/module_next_state[3] , \edb_top_inst/la0/axi_crc_i/n150 , 
        \edb_top_inst/ceg_net221 , \edb_top_inst/la0/axi_crc_i/n149 , \edb_top_inst/la0/axi_crc_i/n148 , 
        \edb_top_inst/la0/axi_crc_i/n147 , \edb_top_inst/la0/axi_crc_i/n146 , 
        \edb_top_inst/la0/axi_crc_i/n145 , \edb_top_inst/la0/axi_crc_i/n144 , 
        \edb_top_inst/la0/axi_crc_i/n143 , \edb_top_inst/la0/axi_crc_i/n142 , 
        \edb_top_inst/la0/axi_crc_i/n141 , \edb_top_inst/la0/axi_crc_i/n140 , 
        \edb_top_inst/la0/axi_crc_i/n139 , \edb_top_inst/la0/axi_crc_i/n138 , 
        \edb_top_inst/la0/axi_crc_i/n137 , \edb_top_inst/la0/axi_crc_i/n136 , 
        \edb_top_inst/la0/axi_crc_i/n135 , \edb_top_inst/la0/axi_crc_i/n134 , 
        \edb_top_inst/la0/axi_crc_i/n133 , \edb_top_inst/la0/axi_crc_i/n132 , 
        \edb_top_inst/la0/axi_crc_i/n131 , \edb_top_inst/la0/axi_crc_i/n130 , 
        \edb_top_inst/la0/axi_crc_i/n129 , \edb_top_inst/la0/axi_crc_i/n128 , 
        \edb_top_inst/la0/axi_crc_i/n127 , \edb_top_inst/la0/axi_crc_i/n126 , 
        \edb_top_inst/la0/axi_crc_i/n125 , \edb_top_inst/la0/axi_crc_i/n124 , 
        \edb_top_inst/la0/axi_crc_i/n123 , \edb_top_inst/la0/axi_crc_i/n122 , 
        \edb_top_inst/la0/axi_crc_i/n121 , \edb_top_inst/la0/axi_crc_i/n120 , 
        \edb_top_inst/la0/axi_crc_i/n119 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n10 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n17 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/equal_9/n3 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n26 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n15 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n9 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n16 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n10 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/equal_9/n3 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n26 , \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n15 , 
        \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n9 , \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/n23 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/genblk1.rise , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/genblk1.fall , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/n18 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n10 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n17 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/equal_9/n3 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n26 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n15 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n9 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n16 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n10 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/equal_9/n3 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n26 , \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n15 , 
        \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n9 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n72 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n38 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n73 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/equal_9/n31 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n82 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n71 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n70 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n69 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n68 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n67 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n66 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n65 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n64 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n63 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n62 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n61 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n60 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n59 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n58 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n57 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n37 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n36 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n35 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n34 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n33 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n32 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n31 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n30 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n29 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n28 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n27 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n26 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n25 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n24 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n23 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n72 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n38 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n73 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/equal_9/n31 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n82 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n71 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n70 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n69 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n68 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n67 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n66 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n65 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n64 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n63 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n62 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n61 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n60 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n59 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n58 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n57 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n37 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n36 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n35 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n34 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n33 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n32 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n31 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n30 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n29 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n28 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n27 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n26 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n25 , \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n24 , 
        \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n40 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n41 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/equal_9/n15 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n50 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n39 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n38 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n37 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n36 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n35 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n34 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n33 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n21 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n20 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n19 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n18 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n17 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n15 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n40 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n41 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/equal_9/n15 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n50 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n39 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n38 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n37 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n36 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n35 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n34 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n33 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n21 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n20 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n19 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n17 , \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n16 , 
        \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n15 , \edb_top_inst/la0/trigger_tu/n47 , 
        \edb_top_inst/la0/genblk2.global_capture_inst/n47 , \edb_top_inst/la0/la_biu_inst/next_state[0] , 
        \edb_top_inst/la0/la_biu_inst/n1182 , \edb_top_inst/la0/la_biu_inst/run_trig_p1 , 
        \edb_top_inst/la0/la_biu_inst/n369 , \edb_top_inst/la0/la_biu_inst/n1285 , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[0] , \edb_top_inst/la0/la_biu_inst/next_fsm_state[0] , 
        \edb_top_inst/ceg_net351 , \edb_top_inst/la0/la_biu_inst/next_state[3] , 
        \edb_top_inst/la0/la_biu_inst/next_state[2] , \edb_top_inst/la0/la_biu_inst/next_state[1] , 
        \edb_top_inst/ceg_net348 , \edb_top_inst/la0/la_biu_inst/fifo_dout[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[2] , \edb_top_inst/la0/la_biu_inst/fifo_dout[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[4] , \edb_top_inst/la0/la_biu_inst/fifo_dout[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[6] , \edb_top_inst/la0/la_biu_inst/fifo_dout[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[8] , \edb_top_inst/la0/la_biu_inst/fifo_dout[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[10] , \edb_top_inst/la0/la_biu_inst/fifo_dout[11] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[12] , \edb_top_inst/la0/la_biu_inst/fifo_dout[13] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[14] , \edb_top_inst/la0/la_biu_inst/fifo_dout[15] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[16] , \edb_top_inst/la0/la_biu_inst/fifo_dout[17] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[18] , \edb_top_inst/la0/la_biu_inst/fifo_dout[19] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[20] , \edb_top_inst/la0/la_biu_inst/fifo_dout[21] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[22] , \edb_top_inst/la0/la_biu_inst/fifo_dout[23] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[24] , \edb_top_inst/la0/la_biu_inst/fifo_dout[25] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[26] , \edb_top_inst/la0/la_biu_inst/fifo_dout[27] , 
        \edb_top_inst/la0/la_biu_inst/fifo_dout[28] , \edb_top_inst/la0/la_biu_inst/fifo_dout[29] , 
        \edb_top_inst/la0/la_biu_inst/next_fsm_state[1] , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data , 
        \edb_top_inst/la0/la_biu_inst/fifo_rstn , \edb_top_inst/la0/la_biu_inst/fifo_pop , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 , \edb_top_inst/la0/la_biu_inst/fifo_push , 
        \edb_top_inst/ceg_net355 , \edb_top_inst/la0/la_biu_inst/n2027 , 
        \edb_top_inst/n341 , \edb_top_inst/n1081 , \edb_top_inst/n1079 , 
        \edb_top_inst/n1077 , \edb_top_inst/n1075 , \edb_top_inst/n1073 , 
        \edb_top_inst/n1071 , \edb_top_inst/n1069 , \edb_top_inst/n1067 , 
        \edb_top_inst/n1066 , \edb_top_inst/n774 , \edb_top_inst/n1064 , 
        \edb_top_inst/n1062 , \edb_top_inst/n1060 , \edb_top_inst/n1058 , 
        \edb_top_inst/n1056 , \edb_top_inst/n1054 , \edb_top_inst/n1052 , 
        \edb_top_inst/n1050 , \edb_top_inst/n1048 , \edb_top_inst/n776 , 
        \edb_top_inst/n1015 , \edb_top_inst/n1013 , \edb_top_inst/n1011 , 
        \edb_top_inst/n1009 , \edb_top_inst/n1007 , \edb_top_inst/n1005 , 
        \edb_top_inst/n1003 , \edb_top_inst/n1001 , \edb_top_inst/n999 , 
        \edb_top_inst/n780 , \edb_top_inst/n956 , \edb_top_inst/n954 , 
        \edb_top_inst/n952 , \edb_top_inst/n950 , \edb_top_inst/n948 , 
        \edb_top_inst/n946 , \edb_top_inst/n944 , \edb_top_inst/n942 , 
        \edb_top_inst/n940 , \edb_top_inst/n939 , \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] , 
        \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] , 
        \edb_top_inst/n778 , \edb_top_inst/n975 , \edb_top_inst/n973 , 
        \edb_top_inst/n971 , \edb_top_inst/n969 , \edb_top_inst/n967 , 
        \edb_top_inst/n965 , \edb_top_inst/n963 , \edb_top_inst/n961 , 
        \edb_top_inst/n959 , \edb_top_inst/n958 , \edb_top_inst/edb_user_dr[65] , 
        \edb_top_inst/edb_user_dr[66] , \edb_top_inst/edb_user_dr[67] , 
        \edb_top_inst/edb_user_dr[68] , \edb_top_inst/edb_user_dr[69] , 
        \edb_top_inst/edb_user_dr[70] , \edb_top_inst/edb_user_dr[71] , 
        \edb_top_inst/edb_user_dr[72] , \edb_top_inst/edb_user_dr[73] , 
        \edb_top_inst/edb_user_dr[74] , \edb_top_inst/edb_user_dr[75] , 
        \edb_top_inst/edb_user_dr[76] , \edb_top_inst/debug_hub_inst/n266 , 
        \edb_top_inst/debug_hub_inst/n95 , \edb_top_inst/edb_user_dr[81] , 
        \edb_top_inst/n941 , \edb_top_inst/n943 , \edb_top_inst/n945 , 
        \edb_top_inst/n947 , \edb_top_inst/n949 , \edb_top_inst/n951 , 
        \edb_top_inst/n953 , \edb_top_inst/n955 , \edb_top_inst/n957 , 
        \edb_top_inst/n960 , \edb_top_inst/n962 , \edb_top_inst/n964 , 
        \edb_top_inst/n966 , \edb_top_inst/n968 , \edb_top_inst/n970 , 
        \edb_top_inst/n972 , \edb_top_inst/n974 , \edb_top_inst/n976 , 
        \edb_top_inst/n1002 , \edb_top_inst/n1004 , \edb_top_inst/n1006 , 
        \edb_top_inst/n1008 , \edb_top_inst/n1010 , \edb_top_inst/n1012 , 
        \edb_top_inst/n1014 , \edb_top_inst/n1016 , \edb_top_inst/n1051 , 
        \edb_top_inst/n1053 , \edb_top_inst/n1055 , \edb_top_inst/n1057 , 
        \edb_top_inst/n1059 , \edb_top_inst/n1061 , \edb_top_inst/n1063 , 
        \edb_top_inst/n1065 , \edb_top_inst/n1068 , \edb_top_inst/n1070 , 
        \edb_top_inst/n1072 , \edb_top_inst/n1074 , \edb_top_inst/n1076 , 
        \edb_top_inst/n1078 , \edb_top_inst/n1080 , \edb_top_inst/n1082 , 
        \edb_top_inst/n1085 , \edb_top_inst/n1087 , \edb_top_inst/n1089 , 
        \edb_top_inst/n1104 , \edb_top_inst/n1106 , \edb_top_inst/n1108 , 
        \edb_top_inst/n1110 , \edb_top_inst/n1112 , \edb_top_inst/n1114 , 
        \edb_top_inst/n1116 , \edb_top_inst/n1118 , \edb_top_inst/n1120 , 
        \edb_top_inst/n1122 , \edb_top_inst/n1124 , \edb_top_inst/n1126 , 
        \edb_top_inst/n1128 , \edb_top_inst/n1130 , \edb_top_inst/n1132 , 
        \edb_top_inst/n1134 , \edb_top_inst/n1136 , \edb_top_inst/n1138 , 
        \edb_top_inst/n1140 , \edb_top_inst/n1142 , \edb_top_inst/n1144 , 
        \edb_top_inst/n1146 , \edb_top_inst/n1148 , \edb_top_inst/n1150 , 
        \edb_top_inst/n1165 , \edb_top_inst/n1167 , \edb_top_inst/n1169 , 
        \edb_top_inst/n1171 , \edb_top_inst/n1173 , \edb_top_inst/n1178 , 
        \edb_top_inst/n1180 , \edb_top_inst/n1182 , \edb_top_inst/n1184 , 
        \edb_top_inst/n2269 , \edb_top_inst/n53 , \edb_top_inst/n1149 , 
        \edb_top_inst/n1147 , \edb_top_inst/n1145 , \edb_top_inst/n1143 , 
        \edb_top_inst/n1141 , \edb_top_inst/n1139 , \edb_top_inst/n1137 , 
        \edb_top_inst/n1135 , \edb_top_inst/n1133 , \edb_top_inst/n1131 , 
        \edb_top_inst/n1129 , \edb_top_inst/n1127 , \edb_top_inst/n1125 , 
        \edb_top_inst/n1123 , \edb_top_inst/n1121 , \edb_top_inst/n1119 , 
        \edb_top_inst/n1183 , \edb_top_inst/n1117 , \edb_top_inst/n1181 , 
        \edb_top_inst/n1115 , \edb_top_inst/n1179 , \edb_top_inst/n1113 , 
        \edb_top_inst/n1177 , \edb_top_inst/n1111 , \edb_top_inst/n1172 , 
        \edb_top_inst/n1109 , \edb_top_inst/n1170 , \edb_top_inst/n1107 , 
        \edb_top_inst/n1168 , \edb_top_inst/n1105 , \edb_top_inst/n1166 , 
        \edb_top_inst/n1103 , \edb_top_inst/n1164 , \edb_top_inst/n1101 , 
        \edb_top_inst/n1162 , \edb_top_inst/n55 , \edb_top_inst/n1088 , 
        \edb_top_inst/n1086 , \edb_top_inst/n1084 , \edb_top_inst/n1083 , 
        \clk~O , \jtag_inst1_TCK~O , n4503, n4504, n4505, n4506, 
        n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, 
        n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, 
        n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, 
        n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, 
        n4540, n4541, n4542, n4543;
    
    EFX_LUT4 LUT__6745 (.I0(\state[1] ), .I1(RX_DV), .O(ceg_net133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__6745.LUTMASK = 16'hbbbb;
    EFX_FF \data[0]~FF  (.D(\received_data[0] ), .CE(ceg_net98), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\data[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \data[0]~FF .CE_POLARITY = 1'b0;
    defparam \data[0]~FF .SR_POLARITY = 1'b1;
    defparam \data[0]~FF .D_POLARITY = 1'b1;
    defparam \data[0]~FF .SR_SYNC = 1'b1;
    defparam \data[0]~FF .SR_VALUE = 1'b0;
    defparam \data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DV~FF  (.D(\state[1] ), .CE(ceg_net127), .CLK(\clk~O ), .SR(1'b0), 
           .Q(DV)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \DV~FF .CLK_POLARITY = 1'b1;
    defparam \DV~FF .CE_POLARITY = 1'b0;
    defparam \DV~FF .SR_POLARITY = 1'b1;
    defparam \DV~FF .D_POLARITY = 1'b0;
    defparam \DV~FF .SR_SYNC = 1'b1;
    defparam \DV~FF .SR_VALUE = 1'b0;
    defparam \DV~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_command~FF  (.D(\state[0] ), .CE(ceg_net130), .CLK(\clk~O ), 
           .SR(1'b0), .Q(led_command)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \led_command~FF .CLK_POLARITY = 1'b1;
    defparam \led_command~FF .CE_POLARITY = 1'b0;
    defparam \led_command~FF .SR_POLARITY = 1'b1;
    defparam \led_command~FF .D_POLARITY = 1'b0;
    defparam \led_command~FF .SR_SYNC = 1'b1;
    defparam \led_command~FF .SR_VALUE = 1'b0;
    defparam \led_command~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \led_data~FF  (.D(n257_2), .CE(ceg_net133), .CLK(\clk~O ), 
           .SR(1'b0), .Q(led_data)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \led_data~FF .CLK_POLARITY = 1'b1;
    defparam \led_data~FF .CE_POLARITY = 1'b0;
    defparam \led_data~FF .SR_POLARITY = 1'b1;
    defparam \led_data~FF .D_POLARITY = 1'b1;
    defparam \led_data~FF .SR_SYNC = 1'b1;
    defparam \led_data~FF .SR_VALUE = 1'b0;
    defparam \led_data~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i[0]~FF  (.D(n62_2), .CE(ceg_net108), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\i[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \i[0]~FF .CLK_POLARITY = 1'b1;
    defparam \i[0]~FF .CE_POLARITY = 1'b0;
    defparam \i[0]~FF .SR_POLARITY = 1'b1;
    defparam \i[0]~FF .D_POLARITY = 1'b1;
    defparam \i[0]~FF .SR_SYNC = 1'b1;
    defparam \i[0]~FF .SR_VALUE = 1'b0;
    defparam \i[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \transmitter_select[0]~FF  (.D(\equal_4/n3 ), .CE(ceg_net120), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\transmitter_select[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \transmitter_select[0]~FF .CLK_POLARITY = 1'b1;
    defparam \transmitter_select[0]~FF .CE_POLARITY = 1'b0;
    defparam \transmitter_select[0]~FF .SR_POLARITY = 1'b1;
    defparam \transmitter_select[0]~FF .D_POLARITY = 1'b0;
    defparam \transmitter_select[0]~FF .SR_SYNC = 1'b1;
    defparam \transmitter_select[0]~FF .SR_VALUE = 1'b0;
    defparam \transmitter_select[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_length[0]~FF  (.D(\received_data[0] ), .CE(ceg_net120), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\data_length[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data_length[0]~FF .CLK_POLARITY = 1'b1;
    defparam \data_length[0]~FF .CE_POLARITY = 1'b0;
    defparam \data_length[0]~FF .SR_POLARITY = 1'b1;
    defparam \data_length[0]~FF .D_POLARITY = 1'b1;
    defparam \data_length[0]~FF .SR_SYNC = 1'b1;
    defparam \data_length[0]~FF .SR_VALUE = 1'b0;
    defparam \data_length[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \state[0]~FF  (.D(\state[0] ), .CE(ceg_net138), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \state[0]~FF .CE_POLARITY = 1'b0;
    defparam \state[0]~FF .SR_POLARITY = 1'b1;
    defparam \state[0]~FF .D_POLARITY = 1'b0;
    defparam \state[0]~FF .SR_SYNC = 1'b1;
    defparam \state[0]~FF .SR_VALUE = 1'b0;
    defparam \state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_Clock_Count[0]~FF  (.D(\uart_rx/n375 ), .CE(ceg_net78), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx/r_Clock_Count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_Clock_Count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[0]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx/r_Clock_Count[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_Clock_Count[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_Clock_Count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \RX_DV~FF  (.D(\uart_rx/n407 ), .CE(ceg_net153), .CLK(\clk~O ), 
           .SR(1'b0), .Q(RX_DV)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \RX_DV~FF .CLK_POLARITY = 1'b1;
    defparam \RX_DV~FF .CE_POLARITY = 1'b0;
    defparam \RX_DV~FF .SR_POLARITY = 1'b1;
    defparam \RX_DV~FF .D_POLARITY = 1'b1;
    defparam \RX_DV~FF .SR_SYNC = 1'b1;
    defparam \RX_DV~FF .SR_VALUE = 1'b0;
    defparam \RX_DV~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_RX_Byte[0]~FF  (.D(rx), .CE(\uart_rx/n444 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\uart_rx/r_RX_Byte[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_RX_Byte[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_RX_Byte[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_RX_Byte[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_Bit_Index[0]~FF  (.D(\uart_rx/n382 ), .CE(ceg_net146), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx/r_Bit_Index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_Bit_Index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_Bit_Index[0]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx/r_Bit_Index[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_Bit_Index[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_Bit_Index[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_Bit_Index[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_Bit_Index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_SM_Main[0]~FF  (.D(\uart_rx/n372 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(\uart_rx/r_SM_Main[2] ), .Q(\uart_rx/r_SM_Main[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_SM_Main[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_SM_Main[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx/r_SM_Main[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_SM_Main[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_SM_Main[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_SM_Main[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_SM_Main[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_Clock_Count[1]~FF  (.D(\uart_rx/n316 ), .CE(ceg_net78), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx/r_Clock_Count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_Clock_Count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[1]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx/r_Clock_Count[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_Clock_Count[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_Clock_Count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_Clock_Count[2]~FF  (.D(\uart_rx/n319 ), .CE(ceg_net78), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx/r_Clock_Count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_Clock_Count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[2]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx/r_Clock_Count[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_Clock_Count[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_Clock_Count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_Clock_Count[3]~FF  (.D(\uart_rx/n322 ), .CE(ceg_net78), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx/r_Clock_Count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_Clock_Count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[3]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx/r_Clock_Count[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[3]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_Clock_Count[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_Clock_Count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_Clock_Count[4]~FF  (.D(\uart_rx/n325 ), .CE(ceg_net78), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx/r_Clock_Count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_Clock_Count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[4]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx/r_Clock_Count[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[4]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_Clock_Count[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_Clock_Count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_Clock_Count[5]~FF  (.D(\uart_rx/n328 ), .CE(ceg_net78), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx/r_Clock_Count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_Clock_Count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[5]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx/r_Clock_Count[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[5]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_Clock_Count[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_Clock_Count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_Clock_Count[6]~FF  (.D(\uart_rx/n331 ), .CE(ceg_net78), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx/r_Clock_Count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_Clock_Count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[6]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx/r_Clock_Count[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[6]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_Clock_Count[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_Clock_Count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_Clock_Count[7]~FF  (.D(\uart_rx/n334 ), .CE(ceg_net78), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx/r_Clock_Count[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_Clock_Count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[7]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx/r_Clock_Count[7]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[7]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_Clock_Count[7]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_Clock_Count[7]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_Clock_Count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_RX_Byte[1]~FF  (.D(rx), .CE(\uart_rx/n429 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\uart_rx/r_RX_Byte[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_RX_Byte[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_RX_Byte[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_RX_Byte[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_RX_Byte[2]~FF  (.D(rx), .CE(\uart_rx/n431 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\uart_rx/r_RX_Byte[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_RX_Byte[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_RX_Byte[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_RX_Byte[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_RX_Byte[3]~FF  (.D(rx), .CE(\uart_rx/n433 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\uart_rx/r_RX_Byte[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_RX_Byte[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[3]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[3]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_RX_Byte[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_RX_Byte[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_RX_Byte[4]~FF  (.D(rx), .CE(\uart_rx/n435 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\uart_rx/r_RX_Byte[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_RX_Byte[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[4]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[4]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_RX_Byte[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_RX_Byte[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_RX_Byte[5]~FF  (.D(rx), .CE(\uart_rx/n437 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\uart_rx/r_RX_Byte[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_RX_Byte[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[5]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[5]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_RX_Byte[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_RX_Byte[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_RX_Byte[6]~FF  (.D(rx), .CE(\uart_rx/n439 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\uart_rx/r_RX_Byte[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_RX_Byte[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[6]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[6]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_RX_Byte[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_RX_Byte[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_RX_Byte[7]~FF  (.D(rx), .CE(\uart_rx/n441 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\uart_rx/r_RX_Byte[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_RX_Byte[7]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[7]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[7]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[7]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_RX_Byte[7]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_RX_Byte[7]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_RX_Byte[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_Bit_Index[1]~FF  (.D(\uart_rx/n359 ), .CE(ceg_net146), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx/r_Bit_Index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_Bit_Index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_Bit_Index[1]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx/r_Bit_Index[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_Bit_Index[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_Bit_Index[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_Bit_Index[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_Bit_Index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_Bit_Index[2]~FF  (.D(\uart_rx/n363 ), .CE(ceg_net146), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_rx/r_Bit_Index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_Bit_Index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_Bit_Index[2]~FF .CE_POLARITY = 1'b0;
    defparam \uart_rx/r_Bit_Index[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_Bit_Index[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_Bit_Index[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_Bit_Index[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_Bit_Index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_SM_Main[1]~FF  (.D(\uart_rx/n309 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(\uart_rx/r_SM_Main[2] ), .Q(\uart_rx/r_SM_Main[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_SM_Main[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_SM_Main[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx/r_SM_Main[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_rx/r_SM_Main[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_rx/r_SM_Main[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_SM_Main[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_SM_Main[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_rx/r_SM_Main[2]~FF  (.D(\uart_rx/n43 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(\uart_rx/n385 ), .Q(\uart_rx/r_SM_Main[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_RX.v(118)
    defparam \uart_rx/r_SM_Main[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_rx/r_SM_Main[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_rx/r_SM_Main[2]~FF .SR_POLARITY = 1'b0;
    defparam \uart_rx/r_SM_Main[2]~FF .D_POLARITY = 1'b0;
    defparam \uart_rx/r_SM_Main[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_rx/r_SM_Main[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_rx/r_SM_Main[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data[1]~FF  (.D(\received_data[1] ), .CE(ceg_net98), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\data[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data[1]~FF .CLK_POLARITY = 1'b1;
    defparam \data[1]~FF .CE_POLARITY = 1'b0;
    defparam \data[1]~FF .SR_POLARITY = 1'b1;
    defparam \data[1]~FF .D_POLARITY = 1'b1;
    defparam \data[1]~FF .SR_SYNC = 1'b1;
    defparam \data[1]~FF .SR_VALUE = 1'b0;
    defparam \data[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data[2]~FF  (.D(\received_data[2] ), .CE(ceg_net98), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\data[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data[2]~FF .CLK_POLARITY = 1'b1;
    defparam \data[2]~FF .CE_POLARITY = 1'b0;
    defparam \data[2]~FF .SR_POLARITY = 1'b1;
    defparam \data[2]~FF .D_POLARITY = 1'b1;
    defparam \data[2]~FF .SR_SYNC = 1'b1;
    defparam \data[2]~FF .SR_VALUE = 1'b0;
    defparam \data[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data[3]~FF  (.D(\received_data[3] ), .CE(ceg_net98), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\data[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data[3]~FF .CLK_POLARITY = 1'b1;
    defparam \data[3]~FF .CE_POLARITY = 1'b0;
    defparam \data[3]~FF .SR_POLARITY = 1'b1;
    defparam \data[3]~FF .D_POLARITY = 1'b1;
    defparam \data[3]~FF .SR_SYNC = 1'b1;
    defparam \data[3]~FF .SR_VALUE = 1'b0;
    defparam \data[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data[4]~FF  (.D(\received_data[4] ), .CE(ceg_net98), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\data[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \data[4]~FF .CE_POLARITY = 1'b0;
    defparam \data[4]~FF .SR_POLARITY = 1'b1;
    defparam \data[4]~FF .D_POLARITY = 1'b1;
    defparam \data[4]~FF .SR_SYNC = 1'b1;
    defparam \data[4]~FF .SR_VALUE = 1'b0;
    defparam \data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data[5]~FF  (.D(\received_data[5] ), .CE(ceg_net98), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\data[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data[5]~FF .CLK_POLARITY = 1'b1;
    defparam \data[5]~FF .CE_POLARITY = 1'b0;
    defparam \data[5]~FF .SR_POLARITY = 1'b1;
    defparam \data[5]~FF .D_POLARITY = 1'b1;
    defparam \data[5]~FF .SR_SYNC = 1'b1;
    defparam \data[5]~FF .SR_VALUE = 1'b0;
    defparam \data[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data[6]~FF  (.D(\received_data[6] ), .CE(ceg_net98), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\data[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data[6]~FF .CLK_POLARITY = 1'b1;
    defparam \data[6]~FF .CE_POLARITY = 1'b0;
    defparam \data[6]~FF .SR_POLARITY = 1'b1;
    defparam \data[6]~FF .D_POLARITY = 1'b1;
    defparam \data[6]~FF .SR_SYNC = 1'b1;
    defparam \data[6]~FF .SR_VALUE = 1'b0;
    defparam \data[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data[7]~FF  (.D(\received_data[7] ), .CE(ceg_net98), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\data[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data[7]~FF .CLK_POLARITY = 1'b1;
    defparam \data[7]~FF .CE_POLARITY = 1'b0;
    defparam \data[7]~FF .SR_POLARITY = 1'b1;
    defparam \data[7]~FF .D_POLARITY = 1'b1;
    defparam \data[7]~FF .SR_SYNC = 1'b1;
    defparam \data[7]~FF .SR_VALUE = 1'b0;
    defparam \data[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i[1]~FF  (.D(n61_2), .CE(ceg_net108), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\i[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \i[1]~FF .CLK_POLARITY = 1'b1;
    defparam \i[1]~FF .CE_POLARITY = 1'b0;
    defparam \i[1]~FF .SR_POLARITY = 1'b1;
    defparam \i[1]~FF .D_POLARITY = 1'b1;
    defparam \i[1]~FF .SR_SYNC = 1'b1;
    defparam \i[1]~FF .SR_VALUE = 1'b0;
    defparam \i[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i[2]~FF  (.D(n60_2), .CE(ceg_net108), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\i[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \i[2]~FF .CLK_POLARITY = 1'b1;
    defparam \i[2]~FF .CE_POLARITY = 1'b0;
    defparam \i[2]~FF .SR_POLARITY = 1'b1;
    defparam \i[2]~FF .D_POLARITY = 1'b1;
    defparam \i[2]~FF .SR_SYNC = 1'b1;
    defparam \i[2]~FF .SR_VALUE = 1'b0;
    defparam \i[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i[3]~FF  (.D(n59_2), .CE(ceg_net108), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\i[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \i[3]~FF .CLK_POLARITY = 1'b1;
    defparam \i[3]~FF .CE_POLARITY = 1'b0;
    defparam \i[3]~FF .SR_POLARITY = 1'b1;
    defparam \i[3]~FF .D_POLARITY = 1'b1;
    defparam \i[3]~FF .SR_SYNC = 1'b1;
    defparam \i[3]~FF .SR_VALUE = 1'b0;
    defparam \i[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i[4]~FF  (.D(n58_2), .CE(ceg_net108), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\i[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \i[4]~FF .CLK_POLARITY = 1'b1;
    defparam \i[4]~FF .CE_POLARITY = 1'b0;
    defparam \i[4]~FF .SR_POLARITY = 1'b1;
    defparam \i[4]~FF .D_POLARITY = 1'b1;
    defparam \i[4]~FF .SR_SYNC = 1'b1;
    defparam \i[4]~FF .SR_VALUE = 1'b0;
    defparam \i[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i[5]~FF  (.D(n57), .CE(ceg_net108), .CLK(\clk~O ), .SR(1'b0), 
           .Q(\i[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \i[5]~FF .CLK_POLARITY = 1'b1;
    defparam \i[5]~FF .CE_POLARITY = 1'b0;
    defparam \i[5]~FF .SR_POLARITY = 1'b1;
    defparam \i[5]~FF .D_POLARITY = 1'b1;
    defparam \i[5]~FF .SR_SYNC = 1'b1;
    defparam \i[5]~FF .SR_VALUE = 1'b0;
    defparam \i[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \transmitter_select[1]~FF  (.D(\equal_5/n3 ), .CE(ceg_net120), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\transmitter_select[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \transmitter_select[1]~FF .CLK_POLARITY = 1'b1;
    defparam \transmitter_select[1]~FF .CE_POLARITY = 1'b0;
    defparam \transmitter_select[1]~FF .SR_POLARITY = 1'b1;
    defparam \transmitter_select[1]~FF .D_POLARITY = 1'b0;
    defparam \transmitter_select[1]~FF .SR_SYNC = 1'b1;
    defparam \transmitter_select[1]~FF .SR_VALUE = 1'b0;
    defparam \transmitter_select[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_length[1]~FF  (.D(\received_data[1] ), .CE(ceg_net120), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\data_length[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data_length[1]~FF .CLK_POLARITY = 1'b1;
    defparam \data_length[1]~FF .CE_POLARITY = 1'b0;
    defparam \data_length[1]~FF .SR_POLARITY = 1'b1;
    defparam \data_length[1]~FF .D_POLARITY = 1'b1;
    defparam \data_length[1]~FF .SR_SYNC = 1'b1;
    defparam \data_length[1]~FF .SR_VALUE = 1'b0;
    defparam \data_length[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_length[2]~FF  (.D(\received_data[2] ), .CE(ceg_net120), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\data_length[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data_length[2]~FF .CLK_POLARITY = 1'b1;
    defparam \data_length[2]~FF .CE_POLARITY = 1'b0;
    defparam \data_length[2]~FF .SR_POLARITY = 1'b1;
    defparam \data_length[2]~FF .D_POLARITY = 1'b1;
    defparam \data_length[2]~FF .SR_SYNC = 1'b1;
    defparam \data_length[2]~FF .SR_VALUE = 1'b0;
    defparam \data_length[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_length[3]~FF  (.D(\received_data[3] ), .CE(ceg_net120), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\data_length[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data_length[3]~FF .CLK_POLARITY = 1'b1;
    defparam \data_length[3]~FF .CE_POLARITY = 1'b0;
    defparam \data_length[3]~FF .SR_POLARITY = 1'b1;
    defparam \data_length[3]~FF .D_POLARITY = 1'b1;
    defparam \data_length[3]~FF .SR_SYNC = 1'b1;
    defparam \data_length[3]~FF .SR_VALUE = 1'b0;
    defparam \data_length[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_length[4]~FF  (.D(\received_data[4] ), .CE(ceg_net120), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\data_length[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data_length[4]~FF .CLK_POLARITY = 1'b1;
    defparam \data_length[4]~FF .CE_POLARITY = 1'b0;
    defparam \data_length[4]~FF .SR_POLARITY = 1'b1;
    defparam \data_length[4]~FF .D_POLARITY = 1'b1;
    defparam \data_length[4]~FF .SR_SYNC = 1'b1;
    defparam \data_length[4]~FF .SR_VALUE = 1'b0;
    defparam \data_length[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_length[5]~FF  (.D(\received_data[5] ), .CE(ceg_net120), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\data_length[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \data_length[5]~FF .CLK_POLARITY = 1'b1;
    defparam \data_length[5]~FF .CE_POLARITY = 1'b0;
    defparam \data_length[5]~FF .SR_POLARITY = 1'b1;
    defparam \data_length[5]~FF .D_POLARITY = 1'b1;
    defparam \data_length[5]~FF .SR_SYNC = 1'b1;
    defparam \data_length[5]~FF .SR_VALUE = 1'b0;
    defparam \data_length[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_Clock_Count[0]~FF  (.D(\uart_tx1/n119 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_Clock_Count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_Clock_Count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_Clock_Count[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_Clock_Count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx1~FF  (.D(\uart_tx1/n110 ), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(tx1)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \tx1~FF .CLK_POLARITY = 1'b1;
    defparam \tx1~FF .CE_POLARITY = 1'b1;
    defparam \tx1~FF .SR_POLARITY = 1'b1;
    defparam \tx1~FF .D_POLARITY = 1'b1;
    defparam \tx1~FF .SR_SYNC = 1'b1;
    defparam \tx1~FF .SR_VALUE = 1'b0;
    defparam \tx1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_Bit_Index[0]~FF  (.D(\uart_tx1/select_38/Select_0/n3 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_Bit_Index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_Bit_Index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_Bit_Index[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_Bit_Index[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_Bit_Index[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_Bit_Index[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_Bit_Index[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_Bit_Index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_TX_Data[0]~FF  (.D(\data_to_transmitter[0] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_TX_Data[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_TX_Data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_TX_Data[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_TX_Data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_SM_Main[0]~FF  (.D(\uart_tx1/n138 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\uart_tx1/r_SM_Main[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_SM_Main[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_SM_Main[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_SM_Main[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_SM_Main[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_SM_Main[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_SM_Main[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_SM_Main[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_Clock_Count[1]~FF  (.D(\uart_tx1/n118 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_Clock_Count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_Clock_Count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_Clock_Count[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_Clock_Count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_Clock_Count[2]~FF  (.D(\uart_tx1/n117 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_Clock_Count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_Clock_Count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_Clock_Count[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_Clock_Count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_Clock_Count[3]~FF  (.D(\uart_tx1/n116 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_Clock_Count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_Clock_Count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[3]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[3]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_Clock_Count[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_Clock_Count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_Clock_Count[4]~FF  (.D(\uart_tx1/n115 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_Clock_Count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_Clock_Count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[4]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[4]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_Clock_Count[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_Clock_Count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_Clock_Count[5]~FF  (.D(\uart_tx1/n114 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_Clock_Count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_Clock_Count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[5]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[5]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_Clock_Count[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_Clock_Count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_Clock_Count[6]~FF  (.D(\uart_tx1/n113 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_Clock_Count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_Clock_Count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[6]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[6]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_Clock_Count[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_Clock_Count[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_Clock_Count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_Bit_Index[1]~FF  (.D(\uart_tx1/n122 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_Bit_Index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_Bit_Index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_Bit_Index[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_Bit_Index[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_Bit_Index[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_Bit_Index[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_Bit_Index[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_Bit_Index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_Bit_Index[2]~FF  (.D(\uart_tx1/n121 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_Bit_Index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_Bit_Index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_Bit_Index[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_Bit_Index[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_Bit_Index[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_Bit_Index[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_Bit_Index[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_Bit_Index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_TX_Data[1]~FF  (.D(\data_to_transmitter[1] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_TX_Data[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_TX_Data[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_TX_Data[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_TX_Data[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_TX_Data[2]~FF  (.D(\data_to_transmitter[2] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_TX_Data[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_TX_Data[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_TX_Data[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_TX_Data[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_TX_Data[3]~FF  (.D(\data_to_transmitter[3] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_TX_Data[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_TX_Data[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[3]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[3]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_TX_Data[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_TX_Data[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_TX_Data[4]~FF  (.D(\data_to_transmitter[4] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_TX_Data[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_TX_Data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[4]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[4]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_TX_Data[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_TX_Data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_TX_Data[5]~FF  (.D(\data_to_transmitter[5] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_TX_Data[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_TX_Data[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[5]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[5]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_TX_Data[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_TX_Data[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_TX_Data[6]~FF  (.D(\data_to_transmitter[6] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_TX_Data[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_TX_Data[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[6]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[6]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_TX_Data[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_TX_Data[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_TX_Data[7]~FF  (.D(\data_to_transmitter[7] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx1/r_TX_Data[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_TX_Data[7]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[7]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[7]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[7]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_TX_Data[7]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_TX_Data[7]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_TX_Data[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx1/r_SM_Main[1]~FF  (.D(\uart_tx1/n137 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\uart_tx1/r_SM_Main[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx1/r_SM_Main[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx1/r_SM_Main[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx1/r_SM_Main[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx1/r_SM_Main[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx1/r_SM_Main[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx1/r_SM_Main[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx1/r_SM_Main[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx2~FF  (.D(\uart_tx2/n110 ), .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), 
           .Q(tx2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \tx2~FF .CLK_POLARITY = 1'b1;
    defparam \tx2~FF .CE_POLARITY = 1'b1;
    defparam \tx2~FF .SR_POLARITY = 1'b1;
    defparam \tx2~FF .D_POLARITY = 1'b1;
    defparam \tx2~FF .SR_SYNC = 1'b1;
    defparam \tx2~FF .SR_VALUE = 1'b0;
    defparam \tx2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx2/r_TX_Data[0]~FF  (.D(\data_to_transmitter[8] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx2/r_TX_Data[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx2/r_TX_Data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[0]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[0]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[0]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[0]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx2/r_TX_Data[0]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx2/r_TX_Data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx2/r_TX_Data[1]~FF  (.D(\data_to_transmitter[9] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx2/r_TX_Data[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx2/r_TX_Data[1]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[1]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[1]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[1]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[1]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx2/r_TX_Data[1]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx2/r_TX_Data[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx2/r_TX_Data[2]~FF  (.D(\data_to_transmitter[10] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx2/r_TX_Data[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx2/r_TX_Data[2]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[2]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[2]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[2]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[2]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx2/r_TX_Data[2]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx2/r_TX_Data[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx2/r_TX_Data[3]~FF  (.D(\data_to_transmitter[11] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx2/r_TX_Data[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx2/r_TX_Data[3]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[3]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[3]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[3]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[3]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx2/r_TX_Data[3]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx2/r_TX_Data[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx2/r_TX_Data[4]~FF  (.D(\data_to_transmitter[12] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx2/r_TX_Data[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx2/r_TX_Data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[4]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[4]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[4]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[4]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx2/r_TX_Data[4]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx2/r_TX_Data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx2/r_TX_Data[5]~FF  (.D(\data_to_transmitter[13] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx2/r_TX_Data[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx2/r_TX_Data[5]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[5]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[5]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[5]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[5]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx2/r_TX_Data[5]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx2/r_TX_Data[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx2/r_TX_Data[6]~FF  (.D(\data_to_transmitter[14] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx2/r_TX_Data[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx2/r_TX_Data[6]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[6]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[6]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[6]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[6]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx2/r_TX_Data[6]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx2/r_TX_Data[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \uart_tx2/r_TX_Data[7]~FF  (.D(\data_to_transmitter[15] ), .CE(\uart_tx1/n338 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\uart_tx2/r_TX_Data[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Documents/Dual_TX_Controll/UART_TX.v(122)
    defparam \uart_tx2/r_TX_Data[7]~FF .CLK_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[7]~FF .CE_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[7]~FF .SR_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[7]~FF .D_POLARITY = 1'b1;
    defparam \uart_tx2/r_TX_Data[7]~FF .SR_SYNC = 1'b1;
    defparam \uart_tx2/r_TX_Data[7]~FF .SR_VALUE = 1'b0;
    defparam \uart_tx2/r_TX_Data[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \state[1]~FF  (.D(n257_2), .CE(ceg_net138), .CLK(\clk~O ), 
           .SR(\state[1] ), .Q(\state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/UART_Controller.v(100)
    defparam \state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \state[1]~FF .CE_POLARITY = 1'b0;
    defparam \state[1]~FF .SR_POLARITY = 1'b1;
    defparam \state[1]~FF .D_POLARITY = 1'b1;
    defparam \state[1]~FF .SR_SYNC = 1'b1;
    defparam \state[1]~FF .SR_VALUE = 1'b0;
    defparam \state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig~FF  (.D(\edb_top_inst/la0/n1334 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_run_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_run_trig_imdt~FF  (.D(\edb_top_inst/la0/n1335 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_run_trig_imdt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_run_trig_imdt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_stop_trig~FF  (.D(\edb_top_inst/la0/n1336 ), 
           .CE(\edb_top_inst/ceg_net5 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_stop_trig )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_stop_trig~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_stop_trig~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[0]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[0]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[0]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_soft_reset_in~FF  (.D(\edb_top_inst/la0/n1959 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_soft_reset_in )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3651)
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_soft_reset_in~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[0]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[0] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3680)
    defparam \edb_top_inst/la0/opcode[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[0]~FF  (.D(\edb_top_inst/la0/n2183 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3689)
    defparam \edb_top_inst/la0/bit_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[0]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[0] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[0]~FF  (.D(\edb_top_inst/la0/n2460 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[0]~FF  (.D(\edb_top_inst/la0/module_next_state[0] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3762)
    defparam \edb_top_inst/la0/module_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn_p1~FF  (.D(1'b1), .CE(1'b1), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_soft_reset_in ), .Q(\edb_top_inst/la0/la_resetn_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4072)
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF  (.D(\state[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_resetn~FF  (.D(\edb_top_inst/la0/la_resetn_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_soft_reset_in ), 
           .Q(\edb_top_inst/la0/la_resetn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4072)
    defparam \edb_top_inst/la0/la_resetn~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_resetn~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n2774 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n2789 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n2987 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n3185 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n3200 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n3398 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF  (.D(RX_DV), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n3611 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n3611 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4022 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF  (.D(\transmitter_select[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4460 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4460 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4475 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4673 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4871 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n4886 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5084 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF  (.D(\data_to_transmitter[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5409 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5820 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF  (.D(\data[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6316 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6331 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6529 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6727 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6742 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n6940 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk2.la_capture_mask[0]~FF  (.D(\edb_top_inst/edb_user_dr[0] ), 
           .CE(\edb_top_inst/la0/n7152 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/genblk2.la_capture_mask[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4349)
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[1]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[0]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[0]~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[0]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_capture_pattern[1]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_capture_pattern[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_capture_pattern[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[16]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[17]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[18]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[19]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[20]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[21]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[22]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[23]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[24]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[25]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[26]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[27]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[28]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[29]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[30]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[31]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[32]~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[33]~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[34]~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[35]~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[36]~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[37]~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[38]~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[39]~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[40]~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[41]~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[42]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[43]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[44]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[45]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[46]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[47]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[48]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[49]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[50]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[51]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[52]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[53]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[54]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[55]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[56]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[57]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[58]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[59]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[60]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[61]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[62]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_mask[63]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1390 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_mask[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3624)
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_mask[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[1]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[2]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[3]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[4]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[5]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[6]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[7]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[8]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[9]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[10]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[11]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[12]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[13]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[14]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[15]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_num_trigger[16]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_num_trigger[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_num_trigger[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[1]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[2]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[3]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_window_depth[4]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/la0/n1907 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_window_depth[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3636)
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_window_depth[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[1]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[1] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[2]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[2] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[3]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[3] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[4]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[4] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[5]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[5] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[6]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[6] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[7]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[7] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[8]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[8] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[9]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[9] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[10]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[10] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[11]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[11] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[12]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[12] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[13]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[13] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[14]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[14] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[15]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[15] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[16]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[16] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[17]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[17] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[18]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[18] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[19]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[19] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[20]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[20] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[21]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[21] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[22]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[22] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[23]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[23] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[24]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[24] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/address_counter[25]~FF  (.D(\edb_top_inst/la0/data_to_addr_counter[25] ), 
           .CE(\edb_top_inst/la0/addr_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/address_counter[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3670)
    defparam \edb_top_inst/la0/address_counter[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/address_counter[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3680)
    defparam \edb_top_inst/la0/opcode[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3680)
    defparam \edb_top_inst/la0/opcode[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/opcode[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/la0/op_reg_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/opcode[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3680)
    defparam \edb_top_inst/la0/opcode[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/opcode[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[1]~FF  (.D(\edb_top_inst/la0/n2182 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3689)
    defparam \edb_top_inst/la0/bit_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[2]~FF  (.D(\edb_top_inst/la0/n2181 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3689)
    defparam \edb_top_inst/la0/bit_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[3]~FF  (.D(\edb_top_inst/la0/n2180 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3689)
    defparam \edb_top_inst/la0/bit_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[4]~FF  (.D(\edb_top_inst/la0/n2179 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3689)
    defparam \edb_top_inst/la0/bit_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/bit_count[5]~FF  (.D(\edb_top_inst/la0/n2178 ), 
           .CE(\edb_top_inst/ceg_net26 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/bit_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3689)
    defparam \edb_top_inst/la0/bit_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/bit_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[1]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[1] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[2]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[2] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[3]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[3] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[4]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[4] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[5]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[5] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[6]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[6] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[7]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[7] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[8]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[8] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[9]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[9] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[10]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[10] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[11]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[11] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[12]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[12] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[13]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[13] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[14]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[14] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/word_count[15]~FF  (.D(\edb_top_inst/la0/data_to_word_counter[15] ), 
           .CE(\edb_top_inst/la0/word_ct_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/word_count[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3707)
    defparam \edb_top_inst/la0/word_count[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/word_count[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[1]~FF  (.D(\edb_top_inst/la0/n2459 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[2]~FF  (.D(\edb_top_inst/la0/n2458 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[3]~FF  (.D(\edb_top_inst/la0/n2457 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[4]~FF  (.D(\edb_top_inst/la0/n2456 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[5]~FF  (.D(\edb_top_inst/la0/n2455 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[6]~FF  (.D(\edb_top_inst/la0/n2454 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[7]~FF  (.D(\edb_top_inst/la0/n2453 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[8]~FF  (.D(\edb_top_inst/la0/n2452 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[9]~FF  (.D(\edb_top_inst/la0/n2451 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[10]~FF  (.D(\edb_top_inst/la0/n2450 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[11]~FF  (.D(\edb_top_inst/la0/n2449 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[12]~FF  (.D(\edb_top_inst/la0/n2448 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[13]~FF  (.D(\edb_top_inst/la0/n2447 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[14]~FF  (.D(\edb_top_inst/la0/n2446 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[15]~FF  (.D(\edb_top_inst/la0/n2445 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[16]~FF  (.D(\edb_top_inst/la0/n2444 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[17]~FF  (.D(\edb_top_inst/la0/n2443 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[18]~FF  (.D(\edb_top_inst/la0/n2442 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[19]~FF  (.D(\edb_top_inst/la0/n2441 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[20]~FF  (.D(\edb_top_inst/la0/n2440 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[21]~FF  (.D(\edb_top_inst/la0/n2439 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[22]~FF  (.D(\edb_top_inst/la0/n2438 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[23]~FF  (.D(\edb_top_inst/la0/n2437 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[24]~FF  (.D(\edb_top_inst/la0/n2436 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[25]~FF  (.D(\edb_top_inst/la0/n2435 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[26]~FF  (.D(\edb_top_inst/la0/n2434 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[27]~FF  (.D(\edb_top_inst/la0/n2433 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[28]~FF  (.D(\edb_top_inst/la0/n2432 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[29]~FF  (.D(\edb_top_inst/la0/n2431 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[30]~FF  (.D(\edb_top_inst/la0/n2430 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[31]~FF  (.D(\edb_top_inst/la0/n2429 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[32]~FF  (.D(\edb_top_inst/la0/n2428 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[33]~FF  (.D(\edb_top_inst/la0/n2427 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[34]~FF  (.D(\edb_top_inst/la0/n2426 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[35]~FF  (.D(\edb_top_inst/la0/n2425 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[36]~FF  (.D(\edb_top_inst/la0/n2424 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[37]~FF  (.D(\edb_top_inst/la0/n2423 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[38]~FF  (.D(\edb_top_inst/la0/n2422 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[39]~FF  (.D(\edb_top_inst/la0/n2421 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[40]~FF  (.D(\edb_top_inst/la0/n2420 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[41]~FF  (.D(\edb_top_inst/la0/n2419 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[42]~FF  (.D(\edb_top_inst/la0/n2418 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[43]~FF  (.D(\edb_top_inst/la0/n2417 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[44]~FF  (.D(\edb_top_inst/la0/n2416 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[45]~FF  (.D(\edb_top_inst/la0/n2415 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[46]~FF  (.D(\edb_top_inst/la0/n2414 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[47]~FF  (.D(\edb_top_inst/la0/n2413 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[48]~FF  (.D(\edb_top_inst/la0/n2412 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[49]~FF  (.D(\edb_top_inst/la0/n2411 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[50]~FF  (.D(\edb_top_inst/la0/n2410 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[51]~FF  (.D(\edb_top_inst/la0/n2409 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[52]~FF  (.D(\edb_top_inst/la0/n2408 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[53]~FF  (.D(\edb_top_inst/la0/n2407 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[54]~FF  (.D(\edb_top_inst/la0/n2406 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[55]~FF  (.D(\edb_top_inst/la0/n2405 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[56]~FF  (.D(\edb_top_inst/la0/n2404 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[57]~FF  (.D(\edb_top_inst/la0/n2403 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[58]~FF  (.D(\edb_top_inst/la0/n2402 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[59]~FF  (.D(\edb_top_inst/la0/n2401 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[60]~FF  (.D(\edb_top_inst/la0/n2400 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[61]~FF  (.D(\edb_top_inst/la0/n2399 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[62]~FF  (.D(\edb_top_inst/la0/n2398 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_out_shift_reg[63]~FF  (.D(\edb_top_inst/la0/n2397 ), 
           .CE(\edb_top_inst/ceg_net14 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/data_out_shift_reg[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3720)
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_out_shift_reg[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[1]~FF  (.D(\edb_top_inst/la0/module_next_state[1] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3762)
    defparam \edb_top_inst/la0/module_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[2]~FF  (.D(\edb_top_inst/la0/module_next_state[2] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3762)
    defparam \edb_top_inst/la0/module_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/module_state[3]~FF  (.D(\edb_top_inst/la0/module_next_state[3] ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/module_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3762)
    defparam \edb_top_inst/la0/module_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/module_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[0]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n150 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[1]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n149 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[2]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n148 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[3]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n147 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[4]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n146 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[5]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n145 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[6]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n144 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[7]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n143 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[8]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n142 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[9]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n141 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[10]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n140 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[11]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n139 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[12]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n138 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[13]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n137 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[14]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n136 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[15]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n135 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[16]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n134 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[17]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n133 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[18]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n132 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[19]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n131 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[20]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n130 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[21]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n129 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[22]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n128 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[23]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n127 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[24]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n126 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[25]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n125 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[26]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n124 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[27]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n123 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[28]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n122 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[29]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n121 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[30]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n120 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/crc_data_out[31]~FF  (.D(\edb_top_inst/la0/axi_crc_i/n119 ), 
           .CE(\edb_top_inst/ceg_net221 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/crc_data_out[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(252)
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/crc_data_out[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1]~FF  (.D(\state[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n2774 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n2774 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n2789 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n2987 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n3185 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n3185 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n3200 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n3398 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n16 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n10 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n17 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/equal_9/n3 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.cap_probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n26 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.cap_probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.cap_probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.cap_probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.cap_probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n15 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n9 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n10 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/equal_9/n3 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n26 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n9 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n3611 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4022 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n4022 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF  (.D(\transmitter_select[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.cap_probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.cap_probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5551)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.cap_probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.cap_probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.cap_probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF  (.D(1'b1), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5490)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5551)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/genblk1.rise ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5551)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/genblk1.fall ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5551)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5551)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5551)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5551)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5490)
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n4460 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4475 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4673 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4871 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n4871 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n4886 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5084 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF  (.D(\data_to_transmitter[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2]~FF  (.D(\data_to_transmitter[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3]~FF  (.D(\data_to_transmitter[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4]~FF  (.D(\data_to_transmitter[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5]~FF  (.D(\data_to_transmitter[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6]~FF  (.D(\data_to_transmitter[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7]~FF  (.D(\data_to_transmitter[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8]~FF  (.D(\data_to_transmitter[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9]~FF  (.D(\data_to_transmitter[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10]~FF  (.D(\data_to_transmitter[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11]~FF  (.D(\data_to_transmitter[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12]~FF  (.D(\data_to_transmitter[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13]~FF  (.D(\data_to_transmitter[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14]~FF  (.D(\data_to_transmitter[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15]~FF  (.D(\data_to_transmitter[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n16 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n10 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n17 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/equal_9/n3 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.cap_probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n26 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.cap_probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.cap_probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.cap_probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.cap_probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n15 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n9 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n10 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/equal_9/n3 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n26 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n9 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5409 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5409 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n5424 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n5622 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5820 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5820 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n5835 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[8]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[9]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[10]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[11]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[12]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[13]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[14]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[15]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/la0/n6033 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF  (.D(\data[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF  (.D(\data[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF  (.D(\data[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF  (.D(\data[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF  (.D(\data[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF  (.D(\data[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF  (.D(\data[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4099)
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n72 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n38 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n73 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/equal_9/n31 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.cap_probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n82 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.cap_probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.cap_probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.cap_probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.cap_probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n71 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n70 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n69 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n68 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n67 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n66 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n65 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n64 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n62 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n61 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n60 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n59 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n58 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n57 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n37 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n36 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n35 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n34 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n33 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n32 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n31 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n30 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n29 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n28 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n27 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n26 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n25 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n24 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n72 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n38 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n73 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/equal_9/n31 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n82 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n71 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n70 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n69 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n68 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n67 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n66 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n65 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n64 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n63 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n62 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n61 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n60 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n59 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n58 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n57 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n37 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n36 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n35 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n33 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n32 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n31 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n30 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n29 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n28 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n27 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n26 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n25 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n24 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6316 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6316 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4191)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6331 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6331 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n6331 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n6331 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n6331 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n6331 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n6331 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4207)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6529 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6529 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n6529 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n6529 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n6529 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n6529 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n6529 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4223)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6727 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6727 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4239)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6742 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6742 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n6742 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n6742 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n6742 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n6742 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n6742 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4255)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n6940 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n6940 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n6940 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n6940 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/la0/n6940 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/la0/n6940 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/la0/n6940 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4271)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk2.la_capture_mask[1]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/la0/n7152 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/genblk2.la_capture_mask[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4349)
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk2.la_capture_mask[2]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/la0/n7152 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/genblk2.la_capture_mask[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4349)
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk2.la_capture_mask[3]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/la0/n7152 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/genblk2.la_capture_mask[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4349)
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk2.la_capture_mask[4]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/la0/n7152 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/genblk2.la_capture_mask[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4349)
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk2.la_capture_mask[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n40 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.cap_probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.cap_probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.cap_probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.cap_probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.cap_probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.cap_probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n39 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n38 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n37 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n36 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n35 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n34 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n33 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n21 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n20 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n19 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n17 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n16 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n15 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n40 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n41 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/equal_9/n15 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n50 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n39 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n38 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n37 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n36 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n35 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n34 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n33 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n21 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n20 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n19 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n17 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n16 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n15 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5602)
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/tu_trigger~FF  (.D(\edb_top_inst/la0/trigger_tu/n47 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/tu_trigger )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5732)
    defparam \edb_top_inst/la0/tu_trigger~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/tu_trigger~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/genblk4.cap_fifo_din_p1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/capture_enable~FF  (.D(\edb_top_inst/la0/genblk2.global_capture_inst/n47 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/capture_enable )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5736)
    defparam \edb_top_inst/la0/capture_enable~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/capture_enable~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/capture_enable~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/capture_enable~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/capture_enable~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/capture_enable~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/capture_enable~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[2]~FF  (.D(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[3]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[4]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[5]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[6]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[7]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[8]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[9]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[10]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[11]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[12]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[13]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[14]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[15]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[16]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[17]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[18]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[19]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[20]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[21]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[22]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[23]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[24]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[25]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[26]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[27]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_cu[28]~FF  (.D(\edb_top_inst/la0/genblk4.cap_fifo_din_p1[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_cu[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4396)
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_cu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[3]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[4]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[7]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[8]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[9]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[10]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[11]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[12]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[13]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[14]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[15]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[16]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[17]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[18]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[19]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[20]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[21]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[22]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[23]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[24]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[25]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[26]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[27]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/cap_fifo_din_tu[28]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_cu[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/cap_fifo_din_tu[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4408)
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/cap_fifo_din_tu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1182 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5218)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5018)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF  (.D(\edb_top_inst/la0/la_run_trig_imdt ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5018)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5018)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n369 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/str_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5239)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5254)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff1 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5254)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5254)
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/str_sync_wbff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5264)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5277)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff1 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5277)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF  (.D(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
           .CE(1'b1), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5277)
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state[0] ), 
           .CE(\edb_top_inst/ceg_net351 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5401)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[3] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1182 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5218)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[2] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1182 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5218)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_state[1] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1182 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/curr_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5218)
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/curr_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF  (.D(\edb_top_inst/la0/la_run_trig ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/run_trig_p1 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5018)
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/run_trig_p1~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/biu_ready~FF  (.D(\edb_top_inst/la0/la_biu_inst/n369 ), 
           .CE(\edb_top_inst/ceg_net348 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/biu_ready )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5289)
    defparam \edb_top_inst/la0/biu_ready~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/biu_ready~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF  (.D(\edb_top_inst/la0/address_counter[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n369 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF  (.D(\edb_top_inst/la0/address_counter[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n369 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF  (.D(\edb_top_inst/la0/address_counter[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n369 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF  (.D(\edb_top_inst/la0/address_counter[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n369 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF  (.D(\edb_top_inst/la0/address_counter[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n369 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF  (.D(\edb_top_inst/la0/address_counter[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n369 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF  (.D(\edb_top_inst/la0/address_counter[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n369 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF  (.D(\edb_top_inst/la0/address_counter[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n369 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF  (.D(\edb_top_inst/la0/address_counter[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n369 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF  (.D(\edb_top_inst/la0/address_counter[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n369 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF  (.D(\edb_top_inst/la0/address_counter[25] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n369 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/la_biu_inst/addr_reg[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5299)
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/addr_reg[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[1] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[2] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[3] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[4] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[5] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[6] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[7] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[8] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[9] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[10] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[11]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[11] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[12]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[12] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[13]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[13] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[14]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[14] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[15]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[15] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[16]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[16] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[17]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[17] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[18]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[18] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[19]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[19] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[20]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[20] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[21]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[21] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[22]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[22] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[23]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[23] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[24]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[24] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[25]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[25] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[26]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[26] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[27]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[27] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[28]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[28] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/data_from_biu[29]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_dout[29] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/n1285 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/data_from_biu[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5308)
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/data_from_biu[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] ), 
           .CE(\edb_top_inst/ceg_net351 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_resetn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(5401)
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/axi_fsm_state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_pop ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[0]~FF  (.D(\edb_top_inst/la0/la_sample_cnt[0] ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_push ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF  (.D(\edb_top_inst/la0/capture_enable ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/n2027 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .D_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF  (.D(\edb_top_inst/n341 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF  (.D(\edb_top_inst/n1081 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF  (.D(\edb_top_inst/n1079 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF  (.D(\edb_top_inst/n1077 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF  (.D(\edb_top_inst/n1075 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF  (.D(\edb_top_inst/n1073 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF  (.D(\edb_top_inst/n1071 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF  (.D(\edb_top_inst/n1069 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF  (.D(\edb_top_inst/n1067 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF  (.D(\edb_top_inst/n1066 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF  (.D(\edb_top_inst/n774 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_pop ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF  (.D(\edb_top_inst/n1064 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_pop ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF  (.D(\edb_top_inst/n1062 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_pop ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF  (.D(\edb_top_inst/n1060 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_pop ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF  (.D(\edb_top_inst/n1058 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_pop ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF  (.D(\edb_top_inst/n1056 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_pop ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF  (.D(\edb_top_inst/n1054 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_pop ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF  (.D(\edb_top_inst/n1052 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_pop ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF  (.D(\edb_top_inst/n1050 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_pop ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF  (.D(\edb_top_inst/n1048 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_pop ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF  (.D(\edb_top_inst/n776 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF  (.D(\edb_top_inst/n1015 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF  (.D(\edb_top_inst/n1013 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF  (.D(\edb_top_inst/n1011 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF  (.D(\edb_top_inst/n1009 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF  (.D(\edb_top_inst/n1007 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF  (.D(\edb_top_inst/n1005 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF  (.D(\edb_top_inst/n1003 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF  (.D(\edb_top_inst/n1001 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF  (.D(\edb_top_inst/n999 ), 
           .CE(\edb_top_inst/la0/la_biu_inst/fifo_push ), .CLK(\clk~O ), 
           .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[1]~FF  (.D(\edb_top_inst/n780 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[2]~FF  (.D(\edb_top_inst/n956 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[3]~FF  (.D(\edb_top_inst/n954 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[4]~FF  (.D(\edb_top_inst/n952 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[5]~FF  (.D(\edb_top_inst/n950 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[6]~FF  (.D(\edb_top_inst/n948 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[7]~FF  (.D(\edb_top_inst/n946 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[8]~FF  (.D(\edb_top_inst/n944 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[9]~FF  (.D(\edb_top_inst/n942 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[10]~FF  (.D(\edb_top_inst/n940 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_sample_cnt[11]~FF  (.D(\edb_top_inst/n939 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
           .Q(\edb_top_inst/la0/la_sample_cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4648)
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_sample_cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[11] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[12] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[13] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[14] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[15] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[16] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[17] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[18] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[19] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[20] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[21] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[22] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[23] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[24] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[25] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[26] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[27] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF  (.D(\edb_top_inst/la0/cap_fifo_din_tu[28] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4717)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF  (.D(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] ), 
           .CE(1'b1), .CLK(\clk~O ), .SR(1'b0), .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4539)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF  (.D(\edb_top_inst/n778 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF  (.D(\edb_top_inst/n975 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF  (.D(\edb_top_inst/n973 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF  (.D(\edb_top_inst/n971 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF  (.D(\edb_top_inst/n969 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF  (.D(\edb_top_inst/n967 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF  (.D(\edb_top_inst/n965 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF  (.D(\edb_top_inst/n963 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF  (.D(\edb_top_inst/n961 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF  (.D(\edb_top_inst/n959 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[11]~FF  (.D(\edb_top_inst/n958 ), 
           .CE(\edb_top_inst/ceg_net355 ), .CLK(\clk~O ), .SR(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 ), 
           .Q(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4634)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[11]~FF .CE_POLARITY = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[11]~FF .SR_SYNC = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[1]~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[2]~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[3]~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[4]~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[5]~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[6]~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[7]~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[8]~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[9]~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[10]~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[11]~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/internal_register_select[12]~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/la0/regsel_ld_en ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/la0/internal_register_select[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3565)
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/internal_register_select[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[1]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[2]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[3]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[4]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[5]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[6]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[7]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[8]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[9]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[10]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_VALUE = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[11]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[12]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[13]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[14]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[15]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/la0/la_trig_pos[16]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/la0/n1306 ), .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), 
           .Q(\edb_top_inst/la0/la_trig_pos[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3614)
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/la0/la_trig_pos[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(323)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[0]~FF  (.D(\edb_top_inst/edb_user_dr[1] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(323)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(323)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n266 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/debug_hub_inst/module_id_reg[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(323)
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/debug_hub_inst/module_id_reg[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[1]~FF  (.D(\edb_top_inst/edb_user_dr[2] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[2]~FF  (.D(\edb_top_inst/edb_user_dr[3] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[3]~FF  (.D(\edb_top_inst/edb_user_dr[4] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[4]~FF  (.D(\edb_top_inst/edb_user_dr[5] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[5]~FF  (.D(\edb_top_inst/edb_user_dr[6] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[6]~FF  (.D(\edb_top_inst/edb_user_dr[7] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[7]~FF  (.D(\edb_top_inst/edb_user_dr[8] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[8]~FF  (.D(\edb_top_inst/edb_user_dr[9] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[9]~FF  (.D(\edb_top_inst/edb_user_dr[10] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[10]~FF  (.D(\edb_top_inst/edb_user_dr[11] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[11]~FF  (.D(\edb_top_inst/edb_user_dr[12] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[12]~FF  (.D(\edb_top_inst/edb_user_dr[13] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[13]~FF  (.D(\edb_top_inst/edb_user_dr[14] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[14]~FF  (.D(\edb_top_inst/edb_user_dr[15] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[15]~FF  (.D(\edb_top_inst/edb_user_dr[16] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[16]~FF  (.D(\edb_top_inst/edb_user_dr[17] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[17]~FF  (.D(\edb_top_inst/edb_user_dr[18] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[18]~FF  (.D(\edb_top_inst/edb_user_dr[19] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[19]~FF  (.D(\edb_top_inst/edb_user_dr[20] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[20]~FF  (.D(\edb_top_inst/edb_user_dr[21] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[21]~FF  (.D(\edb_top_inst/edb_user_dr[22] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[22]~FF  (.D(\edb_top_inst/edb_user_dr[23] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[23]~FF  (.D(\edb_top_inst/edb_user_dr[24] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[24]~FF  (.D(\edb_top_inst/edb_user_dr[25] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[24]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[25]~FF  (.D(\edb_top_inst/edb_user_dr[26] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[25]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[26]~FF  (.D(\edb_top_inst/edb_user_dr[27] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[26]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[27]~FF  (.D(\edb_top_inst/edb_user_dr[28] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[27]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[28]~FF  (.D(\edb_top_inst/edb_user_dr[29] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[28]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[29]~FF  (.D(\edb_top_inst/edb_user_dr[30] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[29]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[30]~FF  (.D(\edb_top_inst/edb_user_dr[31] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[30]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[31]~FF  (.D(\edb_top_inst/edb_user_dr[32] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[31]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[32]~FF  (.D(\edb_top_inst/edb_user_dr[33] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[32]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[33]~FF  (.D(\edb_top_inst/edb_user_dr[34] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[33]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[34]~FF  (.D(\edb_top_inst/edb_user_dr[35] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[34]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[35]~FF  (.D(\edb_top_inst/edb_user_dr[36] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[35]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[36]~FF  (.D(\edb_top_inst/edb_user_dr[37] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[36]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[37]~FF  (.D(\edb_top_inst/edb_user_dr[38] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[37]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[38]~FF  (.D(\edb_top_inst/edb_user_dr[39] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[38]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[39]~FF  (.D(\edb_top_inst/edb_user_dr[40] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[39]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[40]~FF  (.D(\edb_top_inst/edb_user_dr[41] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[40]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[41]~FF  (.D(\edb_top_inst/edb_user_dr[42] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[41]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[42]~FF  (.D(\edb_top_inst/edb_user_dr[43] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[42]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[43]~FF  (.D(\edb_top_inst/edb_user_dr[44] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[43]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[44]~FF  (.D(\edb_top_inst/edb_user_dr[45] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[44]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[45]~FF  (.D(\edb_top_inst/edb_user_dr[46] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[45]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[46]~FF  (.D(\edb_top_inst/edb_user_dr[47] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[46]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[47]~FF  (.D(\edb_top_inst/edb_user_dr[48] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[47]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[48]~FF  (.D(\edb_top_inst/edb_user_dr[49] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[48]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[49]~FF  (.D(\edb_top_inst/edb_user_dr[50] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[49]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[50]~FF  (.D(\edb_top_inst/edb_user_dr[51] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[50]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[51]~FF  (.D(\edb_top_inst/edb_user_dr[52] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[51]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[52]~FF  (.D(\edb_top_inst/edb_user_dr[53] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[52]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[53]~FF  (.D(\edb_top_inst/edb_user_dr[54] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[53]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[54]~FF  (.D(\edb_top_inst/edb_user_dr[55] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[54]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[55]~FF  (.D(\edb_top_inst/edb_user_dr[56] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[55]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[56]~FF  (.D(\edb_top_inst/edb_user_dr[57] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[56]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[57]~FF  (.D(\edb_top_inst/edb_user_dr[58] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[57]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[58]~FF  (.D(\edb_top_inst/edb_user_dr[59] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[58]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[59]~FF  (.D(\edb_top_inst/edb_user_dr[60] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[59]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[60]~FF  (.D(\edb_top_inst/edb_user_dr[61] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[60]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[61]~FF  (.D(\edb_top_inst/edb_user_dr[62] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[61]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[62]~FF  (.D(\edb_top_inst/edb_user_dr[63] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[62]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[63]~FF  (.D(\edb_top_inst/edb_user_dr[64] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[63]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[64]~FF  (.D(\edb_top_inst/edb_user_dr[65] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[64]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[65]~FF  (.D(\edb_top_inst/edb_user_dr[66] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[65]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[66]~FF  (.D(\edb_top_inst/edb_user_dr[67] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[66]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[67]~FF  (.D(\edb_top_inst/edb_user_dr[68] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[67]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[68]~FF  (.D(\edb_top_inst/edb_user_dr[69] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[68]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[69]~FF  (.D(\edb_top_inst/edb_user_dr[70] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[69]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[70]~FF  (.D(\edb_top_inst/edb_user_dr[71] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[70]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[71]~FF  (.D(\edb_top_inst/edb_user_dr[72] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[71]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[72]~FF  (.D(\edb_top_inst/edb_user_dr[73] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[72]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[73]~FF  (.D(\edb_top_inst/edb_user_dr[74] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[73]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[74]~FF  (.D(\edb_top_inst/edb_user_dr[75] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[74]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[75]~FF  (.D(\edb_top_inst/edb_user_dr[76] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[75]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[76]~FF  (.D(\edb_top_inst/edb_user_dr[77] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[76]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[77]~FF  (.D(\edb_top_inst/edb_user_dr[78] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[77]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[78]~FF  (.D(\edb_top_inst/edb_user_dr[79] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[78]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[79]~FF  (.D(\edb_top_inst/edb_user_dr[80] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[79]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[80]~FF  (.D(\edb_top_inst/edb_user_dr[81] ), 
           .CE(\edb_top_inst/debug_hub_inst/n95 ), .CLK(\jtag_inst1_TCK~O ), 
           .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[80]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \edb_top_inst/edb_user_dr[81]~FF  (.D(jtag_inst1_TDI), .CE(\edb_top_inst/debug_hub_inst/n95 ), 
           .CLK(\jtag_inst1_TCK~O ), .SR(jtag_inst1_RESET), .Q(\edb_top_inst/edb_user_dr[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_FF=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(316)
    defparam \edb_top_inst/edb_user_dr[81]~FF .CLK_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .CE_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .D_POLARITY = 1'b1;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_SYNC = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_VALUE = 1'b0;
    defparam \edb_top_inst/edb_user_dr[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_LUT4 \edb_top_inst/LUT__3533  (.I0(\edb_top_inst/la0/crc_data_out[0] ), 
            .I1(\edb_top_inst/edb_user_dr[50] ), .I2(\edb_top_inst/la0/crc_data_out[1] ), 
            .I3(\edb_top_inst/edb_user_dr[51] ), .O(\edb_top_inst/n2270 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3533 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3534  (.I0(\edb_top_inst/la0/crc_data_out[2] ), 
            .I1(\edb_top_inst/edb_user_dr[52] ), .I2(\edb_top_inst/la0/crc_data_out[3] ), 
            .I3(\edb_top_inst/edb_user_dr[53] ), .O(\edb_top_inst/n2271 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3534 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3535  (.I0(\edb_top_inst/la0/crc_data_out[4] ), 
            .I1(\edb_top_inst/edb_user_dr[54] ), .I2(\edb_top_inst/la0/crc_data_out[5] ), 
            .I3(\edb_top_inst/edb_user_dr[55] ), .O(\edb_top_inst/n2272 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3535 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3536  (.I0(\edb_top_inst/n2269 ), .I1(\edb_top_inst/n2270 ), 
            .I2(\edb_top_inst/n2271 ), .I3(\edb_top_inst/n2272 ), .O(\edb_top_inst/n2273 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3536 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3537  (.I0(\edb_top_inst/la0/crc_data_out[12] ), 
            .I1(\edb_top_inst/edb_user_dr[62] ), .I2(\edb_top_inst/la0/crc_data_out[13] ), 
            .I3(\edb_top_inst/edb_user_dr[63] ), .O(\edb_top_inst/n2274 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3537 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3538  (.I0(\edb_top_inst/la0/crc_data_out[7] ), 
            .I1(\edb_top_inst/edb_user_dr[57] ), .I2(\edb_top_inst/la0/crc_data_out[14] ), 
            .I3(\edb_top_inst/edb_user_dr[64] ), .O(\edb_top_inst/n2275 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3538 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3539  (.I0(\edb_top_inst/la0/crc_data_out[8] ), 
            .I1(\edb_top_inst/edb_user_dr[58] ), .I2(\edb_top_inst/la0/crc_data_out[9] ), 
            .I3(\edb_top_inst/edb_user_dr[59] ), .O(\edb_top_inst/n2276 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3539 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3540  (.I0(\edb_top_inst/la0/crc_data_out[10] ), 
            .I1(\edb_top_inst/edb_user_dr[60] ), .I2(\edb_top_inst/la0/crc_data_out[11] ), 
            .I3(\edb_top_inst/edb_user_dr[61] ), .O(\edb_top_inst/n2277 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3540 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3541  (.I0(\edb_top_inst/n2274 ), .I1(\edb_top_inst/n2275 ), 
            .I2(\edb_top_inst/n2276 ), .I3(\edb_top_inst/n2277 ), .O(\edb_top_inst/n2278 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3541 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3542  (.I0(\edb_top_inst/la0/crc_data_out[19] ), 
            .I1(\edb_top_inst/edb_user_dr[69] ), .I2(\edb_top_inst/la0/crc_data_out[20] ), 
            .I3(\edb_top_inst/edb_user_dr[70] ), .O(\edb_top_inst/n2279 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3542 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3543  (.I0(\edb_top_inst/la0/crc_data_out[16] ), 
            .I1(\edb_top_inst/edb_user_dr[66] ), .I2(\edb_top_inst/la0/crc_data_out[23] ), 
            .I3(\edb_top_inst/edb_user_dr[73] ), .O(\edb_top_inst/n2280 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3543 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3544  (.I0(\edb_top_inst/la0/crc_data_out[21] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/la0/crc_data_out[22] ), 
            .I3(\edb_top_inst/edb_user_dr[72] ), .O(\edb_top_inst/n2281 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3544 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3545  (.I0(\edb_top_inst/la0/crc_data_out[17] ), 
            .I1(\edb_top_inst/edb_user_dr[67] ), .I2(\edb_top_inst/la0/crc_data_out[18] ), 
            .I3(\edb_top_inst/edb_user_dr[68] ), .O(\edb_top_inst/n2282 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3545 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3546  (.I0(\edb_top_inst/n2279 ), .I1(\edb_top_inst/n2280 ), 
            .I2(\edb_top_inst/n2281 ), .I3(\edb_top_inst/n2282 ), .O(\edb_top_inst/n2283 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3546 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3547  (.I0(\edb_top_inst/la0/crc_data_out[25] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/la0/crc_data_out[26] ), 
            .I3(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n2284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3547 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3548  (.I0(\edb_top_inst/la0/crc_data_out[24] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/la0/crc_data_out[31] ), 
            .I3(\edb_top_inst/edb_user_dr[81] ), .O(\edb_top_inst/n2285 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3548 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3549  (.I0(\edb_top_inst/la0/crc_data_out[27] ), 
            .I1(\edb_top_inst/edb_user_dr[77] ), .I2(\edb_top_inst/la0/crc_data_out[28] ), 
            .I3(\edb_top_inst/edb_user_dr[78] ), .O(\edb_top_inst/n2286 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3549 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3550  (.I0(\edb_top_inst/la0/crc_data_out[29] ), 
            .I1(\edb_top_inst/edb_user_dr[79] ), .I2(\edb_top_inst/la0/crc_data_out[30] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n2287 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3550 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3551  (.I0(\edb_top_inst/n2284 ), .I1(\edb_top_inst/n2285 ), 
            .I2(\edb_top_inst/n2286 ), .I3(\edb_top_inst/n2287 ), .O(\edb_top_inst/n2288 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3551 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3552  (.I0(\edb_top_inst/n2273 ), .I1(\edb_top_inst/n2278 ), 
            .I2(\edb_top_inst/n2283 ), .I3(\edb_top_inst/n2288 ), .O(\edb_top_inst/n2289 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3552 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3553  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/la0/bit_count[1] ), .I2(\edb_top_inst/la0/bit_count[2] ), 
            .I3(\edb_top_inst/la0/bit_count[3] ), .O(\edb_top_inst/n2290 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3553 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3554  (.I0(\edb_top_inst/la0/bit_count[4] ), 
            .I1(\edb_top_inst/la0/bit_count[5] ), .I2(\edb_top_inst/n2290 ), 
            .O(\edb_top_inst/n2291 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3554 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3555  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n2292 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3555 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3556  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n2293 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3556 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3557  (.I0(\edb_top_inst/n2292 ), .I1(\edb_top_inst/n2291 ), 
            .I2(jtag_inst1_UPDATE), .I3(\edb_top_inst/n2293 ), .O(\edb_top_inst/n2294 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3557 .LUTMASK = 16'h0d00;
    EFX_LUT4 \edb_top_inst/LUT__3558  (.I0(\edb_top_inst/n2294 ), .I1(\edb_top_inst/la0/module_state[3] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2295 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f73, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3558 .LUTMASK = 16'h0f73;
    EFX_LUT4 \edb_top_inst/LUT__3559  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/n2295 ), .O(\edb_top_inst/n2296 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3559 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3560  (.I0(\edb_top_inst/n2289 ), .I1(\edb_top_inst/la0/crc_data_out[0] ), 
            .I2(\edb_top_inst/n2296 ), .O(\edb_top_inst/n2297 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3560 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3561  (.I0(\edb_top_inst/la0/biu_ready ), 
            .I1(\edb_top_inst/la0/data_out_shift_reg[0] ), .I2(\edb_top_inst/n2296 ), 
            .O(\edb_top_inst/n2298 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3561 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3562  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n2299 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3562 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__3563  (.I0(\edb_top_inst/la0/opcode[3] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/n2247 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3563 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3564  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n2244 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3564 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3565  (.I0(\edb_top_inst/n2247 ), .I1(\edb_top_inst/la0/bit_count[5] ), 
            .I2(\edb_top_inst/n2244 ), .I3(\edb_top_inst/la0/bit_count[4] ), 
            .O(\edb_top_inst/n2300 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dfe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3565 .LUTMASK = 16'h3dfe;
    EFX_LUT4 \edb_top_inst/LUT__3566  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[1] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[3] ), .O(\edb_top_inst/n2301 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3566 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__3567  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/la0/bit_count[1] ), .I2(\edb_top_inst/la0/bit_count[2] ), 
            .I3(\edb_top_inst/n2301 ), .O(\edb_top_inst/n2302 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe7f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3567 .LUTMASK = 16'hfe7f;
    EFX_LUT4 \edb_top_inst/LUT__3568  (.I0(\edb_top_inst/la0/opcode[1] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[0] ), .O(\edb_top_inst/n1285 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3568 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3569  (.I0(\edb_top_inst/n2301 ), .I1(\edb_top_inst/n1285 ), 
            .O(\edb_top_inst/n2303 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3569 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3570  (.I0(\edb_top_inst/n2300 ), .I1(\edb_top_inst/n2302 ), 
            .I2(\edb_top_inst/la0/bit_count[3] ), .I3(\edb_top_inst/n2303 ), 
            .O(\edb_top_inst/n2304 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3570 .LUTMASK = 16'h1001;
    EFX_LUT4 \edb_top_inst/LUT__3571  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n2305 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3571 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3572  (.I0(\edb_top_inst/n2304 ), .I1(\edb_top_inst/n2305 ), 
            .O(\edb_top_inst/n2306 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3572 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3573  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n2307 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3573 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3574  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[2] ), 
            .I3(\edb_top_inst/la0/word_count[3] ), .O(\edb_top_inst/n2308 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3574 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3575  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/la0/word_count[6] ), 
            .I3(\edb_top_inst/la0/word_count[7] ), .O(\edb_top_inst/n2309 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3575 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3576  (.I0(\edb_top_inst/la0/word_count[8] ), 
            .I1(\edb_top_inst/la0/word_count[12] ), .I2(\edb_top_inst/la0/word_count[14] ), 
            .I3(\edb_top_inst/la0/word_count[15] ), .O(\edb_top_inst/n2310 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3576 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3577  (.I0(\edb_top_inst/la0/word_count[9] ), 
            .I1(\edb_top_inst/la0/word_count[10] ), .I2(\edb_top_inst/la0/word_count[11] ), 
            .I3(\edb_top_inst/la0/word_count[13] ), .O(\edb_top_inst/n2311 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3577 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3578  (.I0(\edb_top_inst/n2308 ), .I1(\edb_top_inst/n2309 ), 
            .I2(\edb_top_inst/n2310 ), .I3(\edb_top_inst/n2311 ), .O(\edb_top_inst/n2312 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3578 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3579  (.I0(\edb_top_inst/n2307 ), .I1(\edb_top_inst/n2293 ), 
            .I2(\edb_top_inst/n2312 ), .I3(jtag_inst1_UPDATE), .O(\edb_top_inst/n2313 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3579 .LUTMASK = 16'h00f4;
    EFX_LUT4 \edb_top_inst/LUT__3580  (.I0(\edb_top_inst/n2299 ), .I1(\edb_top_inst/n2306 ), 
            .I2(\edb_top_inst/n2293 ), .I3(\edb_top_inst/n2313 ), .O(\edb_top_inst/la0/module_next_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3580 .LUTMASK = 16'hf400;
    EFX_LUT4 \edb_top_inst/LUT__3581  (.I0(\edb_top_inst/n2307 ), .I1(\edb_top_inst/n2312 ), 
            .I2(\edb_top_inst/n2294 ), .O(\edb_top_inst/n2314 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3581 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__3582  (.I0(\edb_top_inst/n2314 ), .I1(\edb_top_inst/la0/module_next_state[3] ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/n2293 ), 
            .O(\edb_top_inst/n2315 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3582 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__3583  (.I0(\edb_top_inst/debug_hub_inst/module_id_reg[1] ), 
            .I1(\edb_top_inst/debug_hub_inst/module_id_reg[2] ), .I2(\edb_top_inst/debug_hub_inst/module_id_reg[3] ), 
            .I3(\edb_top_inst/debug_hub_inst/module_id_reg[0] ), .O(\edb_top_inst/n2316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3583 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3584  (.I0(\edb_top_inst/n2298 ), .I1(\edb_top_inst/n2297 ), 
            .I2(\edb_top_inst/n2315 ), .I3(\edb_top_inst/n2316 ), .O(jtag_inst1_TDO)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3584 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__3585  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[40] ), .O(\edb_top_inst/la0/n1334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3585 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3586  (.I0(\edb_top_inst/edb_user_dr[73] ), 
            .I1(\edb_top_inst/edb_user_dr[74] ), .I2(\edb_top_inst/edb_user_dr[75] ), 
            .I3(\edb_top_inst/edb_user_dr[76] ), .O(\edb_top_inst/n2317 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3586 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3587  (.I0(\edb_top_inst/edb_user_dr[71] ), 
            .I1(\edb_top_inst/n2317 ), .O(\edb_top_inst/n2318 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3587 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3588  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/n2318 ), 
            .O(\edb_top_inst/n2319 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3588 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3589  (.I0(\edb_top_inst/edb_user_dr[67] ), 
            .I1(\edb_top_inst/edb_user_dr[68] ), .I2(\edb_top_inst/edb_user_dr[69] ), 
            .O(\edb_top_inst/n2320 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3589 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3590  (.I0(\edb_top_inst/edb_user_dr[81] ), 
            .I1(jtag_inst1_UPDATE), .I2(\edb_top_inst/n2316 ), .O(\edb_top_inst/n2321 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3590 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3591  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[3] ), .I2(\edb_top_inst/n2307 ), 
            .O(\edb_top_inst/n2322 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3591 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3592  (.I0(\edb_top_inst/edb_user_dr[78] ), 
            .I1(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n2323 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3592 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3593  (.I0(\edb_top_inst/edb_user_dr[77] ), 
            .I1(\edb_top_inst/n2321 ), .I2(\edb_top_inst/n2322 ), .I3(\edb_top_inst/n2323 ), 
            .O(\edb_top_inst/la0/regsel_ld_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3593 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3594  (.I0(\edb_top_inst/edb_user_dr[79] ), 
            .I1(\edb_top_inst/la0/regsel_ld_en ), .O(\edb_top_inst/n2324 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3594 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3595  (.I0(\edb_top_inst/edb_user_dr[66] ), 
            .I1(\edb_top_inst/n2324 ), .O(\edb_top_inst/n2325 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3595 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3596  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n2320 ), 
            .I3(\edb_top_inst/n2325 ), .O(\edb_top_inst/n2326 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3596 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3597  (.I0(\edb_top_inst/n2326 ), .I1(\edb_top_inst/n2319 ), 
            .I2(\edb_top_inst/la0/la_soft_reset_in ), .O(\edb_top_inst/ceg_net5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3597 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3598  (.I0(\edb_top_inst/n2319 ), .I1(\edb_top_inst/n2326 ), 
            .O(\edb_top_inst/la0/n1306 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3598 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3599  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[41] ), .O(\edb_top_inst/la0/n1335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3599 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3600  (.I0(\edb_top_inst/la0/la_soft_reset_in ), 
            .I1(\edb_top_inst/edb_user_dr[42] ), .O(\edb_top_inst/la0/n1336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3600 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3601  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/edb_user_dr[64] ), .I2(\edb_top_inst/n2320 ), 
            .I3(\edb_top_inst/n2325 ), .O(\edb_top_inst/n2327 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3601 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3602  (.I0(\edb_top_inst/n2319 ), .I1(\edb_top_inst/n2327 ), 
            .O(\edb_top_inst/la0/n1390 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3602 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3603  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n2320 ), 
            .I3(\edb_top_inst/n2325 ), .O(\edb_top_inst/n2328 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3603 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3604  (.I0(\edb_top_inst/n2319 ), .I1(\edb_top_inst/n2328 ), 
            .O(\edb_top_inst/la0/n1907 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3604 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3605  (.I0(\edb_top_inst/edb_user_dr[66] ), 
            .I1(\edb_top_inst/n2324 ), .O(\edb_top_inst/n2329 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3605 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3606  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n2320 ), 
            .I3(\edb_top_inst/n2329 ), .O(\edb_top_inst/n2330 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3606 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3607  (.I0(\edb_top_inst/edb_user_dr[63] ), 
            .I1(\edb_top_inst/n2319 ), .I2(\edb_top_inst/n2330 ), .O(\edb_top_inst/la0/n1959 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3607 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__3608  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(\edb_top_inst/la0/address_counter[9] ), .I2(\edb_top_inst/la0/address_counter[10] ), 
            .I3(\edb_top_inst/la0/address_counter[11] ), .O(\edb_top_inst/n2331 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3608 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3609  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/la0/address_counter[12] ), .I2(\edb_top_inst/la0/address_counter[13] ), 
            .I3(\edb_top_inst/la0/address_counter[14] ), .O(\edb_top_inst/n2332 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3609 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3610  (.I0(\edb_top_inst/la0/address_counter[4] ), 
            .I1(\edb_top_inst/la0/address_counter[5] ), .I2(\edb_top_inst/la0/address_counter[6] ), 
            .I3(\edb_top_inst/la0/address_counter[7] ), .O(\edb_top_inst/n2333 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3610 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3611  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/la0/address_counter[1] ), .I2(\edb_top_inst/la0/address_counter[2] ), 
            .O(\edb_top_inst/n2334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3611 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3612  (.I0(\edb_top_inst/n2331 ), .I1(\edb_top_inst/n2332 ), 
            .I2(\edb_top_inst/n2333 ), .I3(\edb_top_inst/n2334 ), .O(\edb_top_inst/n2335 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3612 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3613  (.I0(\edb_top_inst/n2335 ), .I1(\edb_top_inst/n53 ), 
            .I2(\edb_top_inst/edb_user_dr[45] ), .I3(\edb_top_inst/n2322 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3613 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3614  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2336 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3614 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3615  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/module_state[0] ), 
            .O(\edb_top_inst/n2337 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3615 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3616  (.I0(\edb_top_inst/n2337 ), .I1(\edb_top_inst/edb_user_dr[81] ), 
            .I2(\edb_top_inst/n2316 ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n2338 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3616 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__3617  (.I0(\edb_top_inst/n2304 ), .I1(\edb_top_inst/n2312 ), 
            .I2(\edb_top_inst/n2336 ), .I3(\edb_top_inst/n2338 ), .O(\edb_top_inst/n2339 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3617 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__3618  (.I0(\edb_top_inst/n2316 ), .I1(jtag_inst1_CAPTURE), 
            .I2(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n2340 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3618 .LUTMASK = 16'h7070;
    EFX_LUT4 \edb_top_inst/LUT__3619  (.I0(\edb_top_inst/n2340 ), .I1(\edb_top_inst/n2312 ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .O(\edb_top_inst/n2341 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3619 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__3620  (.I0(\edb_top_inst/n2337 ), .I1(\edb_top_inst/n2304 ), 
            .I2(\edb_top_inst/n2312 ), .I3(\edb_top_inst/n2341 ), .O(\edb_top_inst/n2342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3620 .LUTMASK = 16'h7f00;
    EFX_LUT4 \edb_top_inst/LUT__3621  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/n2343 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3621 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3622  (.I0(jtag_inst1_CAPTURE), .I1(\edb_top_inst/n2316 ), 
            .O(\edb_top_inst/n2344 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3622 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3623  (.I0(\edb_top_inst/n2344 ), .I1(\edb_top_inst/n2343 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n2345 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3623 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3624  (.I0(\edb_top_inst/edb_user_dr[77] ), 
            .I1(\edb_top_inst/edb_user_dr[78] ), .I2(\edb_top_inst/edb_user_dr[79] ), 
            .I3(\edb_top_inst/edb_user_dr[80] ), .O(\edb_top_inst/n2346 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe1f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3624 .LUTMASK = 16'hfe1f;
    EFX_LUT4 \edb_top_inst/LUT__3625  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/n2307 ), .O(\edb_top_inst/n2347 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3625 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3626  (.I0(\edb_top_inst/n2346 ), .I1(\edb_top_inst/n2347 ), 
            .I2(\edb_top_inst/n2321 ), .O(\edb_top_inst/n2348 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3626 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3627  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/n2345 ), 
            .I3(\edb_top_inst/n2348 ), .O(\edb_top_inst/n2349 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3627 .LUTMASK = 16'h00bf;
    EFX_LUT4 \edb_top_inst/LUT__3628  (.I0(\edb_top_inst/n2342 ), .I1(\edb_top_inst/n2339 ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .I3(\edb_top_inst/n2349 ), 
            .O(\edb_top_inst/n2350 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3628 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__3629  (.I0(\edb_top_inst/n2350 ), .I1(\edb_top_inst/n2322 ), 
            .O(\edb_top_inst/la0/op_reg_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3629 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3630  (.I0(\edb_top_inst/la0/word_count[1] ), 
            .I1(\edb_top_inst/la0/word_count[2] ), .I2(\edb_top_inst/la0/word_count[3] ), 
            .O(\edb_top_inst/n2351 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3630 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__3631  (.I0(\edb_top_inst/n2310 ), .I1(\edb_top_inst/n2311 ), 
            .I2(\edb_top_inst/n2351 ), .I3(\edb_top_inst/n2309 ), .O(\edb_top_inst/n2352 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3631 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3632  (.I0(\edb_top_inst/n2352 ), .I1(\edb_top_inst/la0/module_state[1] ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/n2304 ), 
            .O(\edb_top_inst/n2353 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3632 .LUTMASK = 16'hc100;
    EFX_LUT4 \edb_top_inst/LUT__3633  (.I0(\edb_top_inst/n2307 ), .I1(\edb_top_inst/la0/module_state[3] ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .O(\edb_top_inst/n2354 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3633 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__3634  (.I0(\edb_top_inst/la0/module_state[2] ), 
            .I1(\edb_top_inst/la0/module_state[1] ), .I2(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n2355 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3634 .LUTMASK = 16'h0707;
    EFX_LUT4 \edb_top_inst/LUT__3635  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/biu_ready ), .I2(\edb_top_inst/n2336 ), 
            .I3(\edb_top_inst/n2355 ), .O(\edb_top_inst/n2356 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3635 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__3636  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .O(\edb_top_inst/n2357 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3636 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3637  (.I0(\edb_top_inst/n2312 ), .I1(\edb_top_inst/n2357 ), 
            .O(\edb_top_inst/n2358 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3637 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3638  (.I0(\edb_top_inst/n2356 ), .I1(\edb_top_inst/n2352 ), 
            .I2(\edb_top_inst/n2358 ), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n2359 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3638 .LUTMASK = 16'h000d;
    EFX_LUT4 \edb_top_inst/LUT__3639  (.I0(\edb_top_inst/n2359 ), .I1(\edb_top_inst/n2353 ), 
            .I2(\edb_top_inst/n2354 ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n2360 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fab, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3639 .LUTMASK = 16'h0fab;
    EFX_LUT4 \edb_top_inst/LUT__3640  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n2360 ), .O(\edb_top_inst/la0/addr_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3640 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3641  (.I0(\edb_top_inst/n2299 ), .I1(\edb_top_inst/n2306 ), 
            .I2(\edb_top_inst/n2356 ), .O(\edb_top_inst/n2361 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3641 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__3642  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n2350 ), .I2(\edb_top_inst/n2347 ), .I3(\edb_top_inst/n2361 ), 
            .O(\edb_top_inst/n2362 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3642 .LUTMASK = 16'h4f00;
    EFX_LUT4 \edb_top_inst/LUT__3643  (.I0(\edb_top_inst/la0/bit_count[0] ), 
            .I1(\edb_top_inst/n2362 ), .O(\edb_top_inst/la0/n2183 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3643 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3644  (.I0(\edb_top_inst/n2350 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/n2305 ), 
            .O(\edb_top_inst/n2363 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd300, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3644 .LUTMASK = 16'hd300;
    EFX_LUT4 \edb_top_inst/LUT__3645  (.I0(\edb_top_inst/n2292 ), .I1(\edb_top_inst/n2293 ), 
            .I2(\edb_top_inst/n2363 ), .I3(\edb_top_inst/n2362 ), .O(\edb_top_inst/ceg_net26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3645 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__3646  (.I0(\edb_top_inst/edb_user_dr[29] ), 
            .I1(\edb_top_inst/la0/word_count[0] ), .I2(\edb_top_inst/n2322 ), 
            .O(\edb_top_inst/la0/data_to_word_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3646 .LUTMASK = 16'ha3a3;
    EFX_LUT4 \edb_top_inst/LUT__3647  (.I0(\edb_top_inst/n2350 ), .I1(\edb_top_inst/la0/module_state[0] ), 
            .I2(\edb_top_inst/n2305 ), .I3(\edb_top_inst/n2362 ), .O(\edb_top_inst/la0/word_ct_en )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h10ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3647 .LUTMASK = 16'h10ff;
    EFX_LUT4 \edb_top_inst/LUT__3648  (.I0(\edb_top_inst/la0/internal_register_select[10] ), 
            .I1(\edb_top_inst/la0/internal_register_select[11] ), .O(\edb_top_inst/n2364 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3648 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3649  (.I0(\edb_top_inst/la0/internal_register_select[6] ), 
            .I1(\edb_top_inst/la0/internal_register_select[7] ), .I2(\edb_top_inst/la0/internal_register_select[8] ), 
            .I3(\edb_top_inst/la0/internal_register_select[9] ), .O(\edb_top_inst/n2365 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3649 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3650  (.I0(\edb_top_inst/la0/internal_register_select[1] ), 
            .I1(\edb_top_inst/la0/internal_register_select[2] ), .I2(\edb_top_inst/la0/internal_register_select[4] ), 
            .I3(\edb_top_inst/la0/internal_register_select[5] ), .O(\edb_top_inst/n2366 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3650 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__3651  (.I0(\edb_top_inst/la0/internal_register_select[12] ), 
            .I1(\edb_top_inst/n2364 ), .I2(\edb_top_inst/n2365 ), .I3(\edb_top_inst/n2366 ), 
            .O(\edb_top_inst/n2367 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3651 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3652  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/internal_register_select[0] ), .I2(\edb_top_inst/n2367 ), 
            .O(\edb_top_inst/n2368 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3652 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3653  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/n2367 ), 
            .O(\edb_top_inst/n2369 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3653 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3654  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n2370 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h13f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3654 .LUTMASK = 16'h13f8;
    EFX_LUT4 \edb_top_inst/LUT__3655  (.I0(\edb_top_inst/n2368 ), .I1(\edb_top_inst/la0/la_trig_mask[0] ), 
            .I2(\edb_top_inst/n2370 ), .I3(\edb_top_inst/n2369 ), .O(\edb_top_inst/n2371 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f77, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3655 .LUTMASK = 16'h0f77;
    EFX_LUT4 \edb_top_inst/LUT__3656  (.I0(\edb_top_inst/n2307 ), .I1(\edb_top_inst/n2304 ), 
            .I2(\edb_top_inst/n2305 ), .I3(\edb_top_inst/n2356 ), .O(\edb_top_inst/n2372 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3656 .LUTMASK = 16'h007f;
    EFX_LUT4 \edb_top_inst/LUT__3657  (.I0(\edb_top_inst/la0/data_from_biu[0] ), 
            .I1(\edb_top_inst/n2371 ), .I2(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2373 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3657 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__3658  (.I0(\edb_top_inst/n2344 ), .I1(\edb_top_inst/n2307 ), 
            .I2(\edb_top_inst/la0/module_state[2] ), .I3(\edb_top_inst/n2356 ), 
            .O(\edb_top_inst/n2374 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3037, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3658 .LUTMASK = 16'h3037;
    EFX_LUT4 \edb_top_inst/LUT__3659  (.I0(\edb_top_inst/n2304 ), .I1(\edb_top_inst/la0/module_state[2] ), 
            .I2(\edb_top_inst/n2374 ), .I3(\edb_top_inst/la0/module_state[3] ), 
            .O(\edb_top_inst/n2375 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3659 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__3660  (.I0(\edb_top_inst/la0/data_out_shift_reg[1] ), 
            .I1(\edb_top_inst/n2373 ), .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3660 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3661  (.I0(jtag_inst1_SHIFT), .I1(jtag_inst1_CAPTURE), 
            .I2(\edb_top_inst/n2316 ), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n2376 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3661 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__3662  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n2376 ), .I2(\edb_top_inst/n2307 ), .I3(\edb_top_inst/n2356 ), 
            .O(\edb_top_inst/ceg_net14 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3662 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__3663  (.I0(\edb_top_inst/la0/module_state[3] ), 
            .I1(\edb_top_inst/n2350 ), .I2(\edb_top_inst/n2314 ), .O(\edb_top_inst/la0/module_next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf1f1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3663 .LUTMASK = 16'hf1f1;
    EFX_LUT4 \edb_top_inst/LUT__3664  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .I3(\edb_top_inst/n2317 ), .O(\edb_top_inst/n2377 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3664 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3665  (.I0(\edb_top_inst/n2326 ), .I1(\edb_top_inst/n2377 ), 
            .O(\edb_top_inst/la0/n2774 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3665 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3666  (.I0(\edb_top_inst/n2327 ), .I1(\edb_top_inst/n2377 ), 
            .O(\edb_top_inst/la0/n2789 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3666 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3667  (.I0(\edb_top_inst/edb_user_dr[64] ), 
            .I1(\edb_top_inst/edb_user_dr[65] ), .I2(\edb_top_inst/n2320 ), 
            .I3(\edb_top_inst/n2325 ), .O(\edb_top_inst/n2378 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3667 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3668  (.I0(\edb_top_inst/n2377 ), .I1(\edb_top_inst/n2378 ), 
            .O(\edb_top_inst/la0/n2987 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3668 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3669  (.I0(\edb_top_inst/n2328 ), .I1(\edb_top_inst/n2377 ), 
            .O(\edb_top_inst/la0/n3185 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3669 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3670  (.I0(\edb_top_inst/n2330 ), .I1(\edb_top_inst/n2377 ), 
            .O(\edb_top_inst/la0/n3200 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3670 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3671  (.I0(\edb_top_inst/edb_user_dr[65] ), 
            .I1(\edb_top_inst/edb_user_dr[64] ), .I2(\edb_top_inst/n2320 ), 
            .I3(\edb_top_inst/n2329 ), .O(\edb_top_inst/n2379 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3671 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3672  (.I0(\edb_top_inst/n2377 ), .I1(\edb_top_inst/n2379 ), 
            .O(\edb_top_inst/la0/n3398 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3672 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3673  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/n2318 ), 
            .I3(\edb_top_inst/n2326 ), .O(\edb_top_inst/la0/n3611 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3673 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3674  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/n2318 ), 
            .I3(\edb_top_inst/n2328 ), .O(\edb_top_inst/la0/n4022 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3674 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3675  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .I3(\edb_top_inst/n2317 ), .O(\edb_top_inst/n2380 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3675 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3676  (.I0(\edb_top_inst/n2326 ), .I1(\edb_top_inst/n2380 ), 
            .O(\edb_top_inst/la0/n4460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3676 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3677  (.I0(\edb_top_inst/n2327 ), .I1(\edb_top_inst/n2380 ), 
            .O(\edb_top_inst/la0/n4475 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3677 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3678  (.I0(\edb_top_inst/n2378 ), .I1(\edb_top_inst/n2380 ), 
            .O(\edb_top_inst/la0/n4673 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3678 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3679  (.I0(\edb_top_inst/n2328 ), .I1(\edb_top_inst/n2380 ), 
            .O(\edb_top_inst/la0/n4871 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3679 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3680  (.I0(\edb_top_inst/n2330 ), .I1(\edb_top_inst/n2380 ), 
            .O(\edb_top_inst/la0/n4886 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3680 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3681  (.I0(\edb_top_inst/n2379 ), .I1(\edb_top_inst/n2380 ), 
            .O(\edb_top_inst/la0/n5084 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3681 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3682  (.I0(\edb_top_inst/edb_user_dr[74] ), 
            .I1(\edb_top_inst/edb_user_dr[75] ), .I2(\edb_top_inst/edb_user_dr[76] ), 
            .I3(\edb_top_inst/edb_user_dr[73] ), .O(\edb_top_inst/n2381 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3682 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3683  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[71] ), .I2(\edb_top_inst/edb_user_dr[72] ), 
            .I3(\edb_top_inst/n2381 ), .O(\edb_top_inst/n2382 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3683 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3684  (.I0(\edb_top_inst/n2326 ), .I1(\edb_top_inst/n2382 ), 
            .O(\edb_top_inst/la0/n5409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3684 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3685  (.I0(\edb_top_inst/n2327 ), .I1(\edb_top_inst/n2382 ), 
            .O(\edb_top_inst/la0/n5424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3685 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3686  (.I0(\edb_top_inst/n2378 ), .I1(\edb_top_inst/n2382 ), 
            .O(\edb_top_inst/la0/n5622 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3686 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3687  (.I0(\edb_top_inst/n2328 ), .I1(\edb_top_inst/n2382 ), 
            .O(\edb_top_inst/la0/n5820 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3687 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3688  (.I0(\edb_top_inst/n2330 ), .I1(\edb_top_inst/n2382 ), 
            .O(\edb_top_inst/la0/n5835 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3688 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3689  (.I0(\edb_top_inst/n2379 ), .I1(\edb_top_inst/n2382 ), 
            .O(\edb_top_inst/la0/n6033 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3689 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3690  (.I0(\edb_top_inst/edb_user_dr[70] ), 
            .I1(\edb_top_inst/edb_user_dr[72] ), .I2(\edb_top_inst/edb_user_dr[71] ), 
            .I3(\edb_top_inst/n2381 ), .O(\edb_top_inst/n2383 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3690 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3691  (.I0(\edb_top_inst/n2326 ), .I1(\edb_top_inst/n2383 ), 
            .O(\edb_top_inst/la0/n6316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3691 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3692  (.I0(\edb_top_inst/n2327 ), .I1(\edb_top_inst/n2383 ), 
            .O(\edb_top_inst/la0/n6331 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3692 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3693  (.I0(\edb_top_inst/n2378 ), .I1(\edb_top_inst/n2383 ), 
            .O(\edb_top_inst/la0/n6529 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3693 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3694  (.I0(\edb_top_inst/n2328 ), .I1(\edb_top_inst/n2383 ), 
            .O(\edb_top_inst/la0/n6727 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3694 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3695  (.I0(\edb_top_inst/n2330 ), .I1(\edb_top_inst/n2383 ), 
            .O(\edb_top_inst/la0/n6742 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3695 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3696  (.I0(\edb_top_inst/n2379 ), .I1(\edb_top_inst/n2383 ), 
            .O(\edb_top_inst/la0/n6940 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3696 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3697  (.I0(\edb_top_inst/n2319 ), .I1(\edb_top_inst/n2378 ), 
            .O(\edb_top_inst/la0/n7152 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3697 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3698  (.I0(\edb_top_inst/n2335 ), .I1(\edb_top_inst/n1149 ), 
            .I2(\edb_top_inst/edb_user_dr[46] ), .I3(\edb_top_inst/n2322 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3698 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3699  (.I0(\edb_top_inst/n2335 ), .I1(\edb_top_inst/n1147 ), 
            .I2(\edb_top_inst/edb_user_dr[47] ), .I3(\edb_top_inst/n2322 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3699 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3700  (.I0(\edb_top_inst/n2335 ), .I1(\edb_top_inst/n1145 ), 
            .I2(\edb_top_inst/edb_user_dr[48] ), .I3(\edb_top_inst/n2322 ), 
            .O(\edb_top_inst/la0/data_to_addr_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3700 .LUTMASK = 16'hf044;
    EFX_LUT4 \edb_top_inst/LUT__3701  (.I0(\edb_top_inst/edb_user_dr[49] ), 
            .I1(\edb_top_inst/n1143 ), .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3701 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3702  (.I0(\edb_top_inst/edb_user_dr[50] ), 
            .I1(\edb_top_inst/n1141 ), .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3702 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3703  (.I0(\edb_top_inst/edb_user_dr[51] ), 
            .I1(\edb_top_inst/n1139 ), .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3703 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3704  (.I0(\edb_top_inst/edb_user_dr[52] ), 
            .I1(\edb_top_inst/n1137 ), .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3704 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3705  (.I0(\edb_top_inst/edb_user_dr[53] ), 
            .I1(\edb_top_inst/n1135 ), .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3705 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3706  (.I0(\edb_top_inst/edb_user_dr[54] ), 
            .I1(\edb_top_inst/n1133 ), .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3706 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3707  (.I0(\edb_top_inst/edb_user_dr[55] ), 
            .I1(\edb_top_inst/n1131 ), .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3707 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3708  (.I0(\edb_top_inst/edb_user_dr[56] ), 
            .I1(\edb_top_inst/n1129 ), .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3708 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3709  (.I0(\edb_top_inst/edb_user_dr[57] ), 
            .I1(\edb_top_inst/n1127 ), .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3709 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3710  (.I0(\edb_top_inst/edb_user_dr[58] ), 
            .I1(\edb_top_inst/n1125 ), .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3710 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3711  (.I0(\edb_top_inst/edb_user_dr[59] ), 
            .I1(\edb_top_inst/n1123 ), .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3711 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3712  (.I0(\edb_top_inst/n1121 ), .I1(\edb_top_inst/la0/address_counter[15] ), 
            .I2(\edb_top_inst/n2335 ), .O(\edb_top_inst/n2384 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3712 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__3713  (.I0(\edb_top_inst/n2384 ), .I1(\edb_top_inst/edb_user_dr[60] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3713 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3714  (.I0(\edb_top_inst/n1183 ), .I1(\edb_top_inst/n1119 ), 
            .I2(\edb_top_inst/n2335 ), .O(\edb_top_inst/n2385 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3714 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3715  (.I0(\edb_top_inst/n2385 ), .I1(\edb_top_inst/edb_user_dr[61] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3715 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3716  (.I0(\edb_top_inst/n1181 ), .I1(\edb_top_inst/n1117 ), 
            .I2(\edb_top_inst/n2335 ), .O(\edb_top_inst/n2386 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3716 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3717  (.I0(\edb_top_inst/n2386 ), .I1(\edb_top_inst/edb_user_dr[62] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3717 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3718  (.I0(\edb_top_inst/n1179 ), .I1(\edb_top_inst/n1115 ), 
            .I2(\edb_top_inst/n2335 ), .O(\edb_top_inst/n2387 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3718 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3719  (.I0(\edb_top_inst/n2387 ), .I1(\edb_top_inst/edb_user_dr[63] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3719 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3720  (.I0(\edb_top_inst/n1177 ), .I1(\edb_top_inst/n1113 ), 
            .I2(\edb_top_inst/n2335 ), .O(\edb_top_inst/n2388 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3720 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3721  (.I0(\edb_top_inst/n2388 ), .I1(\edb_top_inst/edb_user_dr[64] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3721 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3722  (.I0(\edb_top_inst/n1172 ), .I1(\edb_top_inst/n1111 ), 
            .I2(\edb_top_inst/n2335 ), .O(\edb_top_inst/n2389 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3722 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3723  (.I0(\edb_top_inst/n2389 ), .I1(\edb_top_inst/edb_user_dr[65] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3723 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3724  (.I0(\edb_top_inst/n1170 ), .I1(\edb_top_inst/n1109 ), 
            .I2(\edb_top_inst/n2335 ), .O(\edb_top_inst/n2390 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3724 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3725  (.I0(\edb_top_inst/n2390 ), .I1(\edb_top_inst/edb_user_dr[66] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3725 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3726  (.I0(\edb_top_inst/n1168 ), .I1(\edb_top_inst/n1107 ), 
            .I2(\edb_top_inst/n2335 ), .O(\edb_top_inst/n2391 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3726 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3727  (.I0(\edb_top_inst/n2391 ), .I1(\edb_top_inst/edb_user_dr[67] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3727 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3728  (.I0(\edb_top_inst/n1166 ), .I1(\edb_top_inst/n1105 ), 
            .I2(\edb_top_inst/n2335 ), .O(\edb_top_inst/n2392 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3728 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3729  (.I0(\edb_top_inst/n2392 ), .I1(\edb_top_inst/edb_user_dr[68] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3729 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3730  (.I0(\edb_top_inst/n1164 ), .I1(\edb_top_inst/n1103 ), 
            .I2(\edb_top_inst/n2335 ), .O(\edb_top_inst/n2393 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3730 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3731  (.I0(\edb_top_inst/n2393 ), .I1(\edb_top_inst/edb_user_dr[69] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3731 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3732  (.I0(\edb_top_inst/n1162 ), .I1(\edb_top_inst/n1101 ), 
            .I2(\edb_top_inst/n2335 ), .O(\edb_top_inst/n2394 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3732 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3733  (.I0(\edb_top_inst/n2394 ), .I1(\edb_top_inst/edb_user_dr[70] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_addr_counter[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3733 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3746  (.I0(\edb_top_inst/n55 ), .I1(\edb_top_inst/n2362 ), 
            .O(\edb_top_inst/la0/n2182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3746 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3747  (.I0(\edb_top_inst/n1088 ), .I1(\edb_top_inst/n2362 ), 
            .O(\edb_top_inst/la0/n2181 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3747 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3748  (.I0(\edb_top_inst/n1086 ), .I1(\edb_top_inst/n2362 ), 
            .O(\edb_top_inst/la0/n2180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3748 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3749  (.I0(\edb_top_inst/n1084 ), .I1(\edb_top_inst/n2362 ), 
            .O(\edb_top_inst/la0/n2179 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3749 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3750  (.I0(\edb_top_inst/n1083 ), .I1(\edb_top_inst/n2362 ), 
            .O(\edb_top_inst/la0/n2178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3750 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3751  (.I0(\edb_top_inst/edb_user_dr[30] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .I2(\edb_top_inst/la0/word_count[0] ), 
            .I3(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haac3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3751 .LUTMASK = 16'haac3;
    EFX_LUT4 \edb_top_inst/LUT__3752  (.I0(\edb_top_inst/la0/word_count[0] ), 
            .I1(\edb_top_inst/la0/word_count[1] ), .O(\edb_top_inst/n2401 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3752 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3753  (.I0(\edb_top_inst/edb_user_dr[31] ), 
            .I1(\edb_top_inst/la0/word_count[2] ), .I2(\edb_top_inst/n2401 ), 
            .I3(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3753 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3754  (.I0(\edb_top_inst/la0/word_count[2] ), 
            .I1(\edb_top_inst/n2401 ), .I2(\edb_top_inst/la0/word_count[3] ), 
            .O(\edb_top_inst/n2402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3754 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__3755  (.I0(\edb_top_inst/n2402 ), .I1(\edb_top_inst/edb_user_dr[32] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3755 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3756  (.I0(\edb_top_inst/edb_user_dr[33] ), 
            .I1(\edb_top_inst/la0/word_count[4] ), .I2(\edb_top_inst/n2308 ), 
            .I3(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3756 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3757  (.I0(\edb_top_inst/la0/word_count[4] ), 
            .I1(\edb_top_inst/n2308 ), .O(\edb_top_inst/n2403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3757 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3758  (.I0(\edb_top_inst/edb_user_dr[34] ), 
            .I1(\edb_top_inst/la0/word_count[5] ), .I2(\edb_top_inst/n2403 ), 
            .I3(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3758 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3759  (.I0(\edb_top_inst/la0/word_count[5] ), 
            .I1(\edb_top_inst/n2403 ), .O(\edb_top_inst/n2404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3759 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3760  (.I0(\edb_top_inst/edb_user_dr[35] ), 
            .I1(\edb_top_inst/la0/word_count[6] ), .I2(\edb_top_inst/n2404 ), 
            .I3(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3760 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3761  (.I0(\edb_top_inst/la0/word_count[6] ), 
            .I1(\edb_top_inst/n2404 ), .O(\edb_top_inst/n2405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3761 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3762  (.I0(\edb_top_inst/edb_user_dr[36] ), 
            .I1(\edb_top_inst/la0/word_count[7] ), .I2(\edb_top_inst/n2405 ), 
            .I3(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3762 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3763  (.I0(\edb_top_inst/n2308 ), .I1(\edb_top_inst/n2309 ), 
            .O(\edb_top_inst/n2406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3763 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3764  (.I0(\edb_top_inst/edb_user_dr[37] ), 
            .I1(\edb_top_inst/la0/word_count[8] ), .I2(\edb_top_inst/n2406 ), 
            .I3(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3764 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3765  (.I0(\edb_top_inst/la0/word_count[8] ), 
            .I1(\edb_top_inst/n2406 ), .I2(\edb_top_inst/la0/word_count[9] ), 
            .O(\edb_top_inst/n2407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3765 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__3766  (.I0(\edb_top_inst/n2407 ), .I1(\edb_top_inst/edb_user_dr[38] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3766 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3767  (.I0(\edb_top_inst/la0/word_count[8] ), 
            .I1(\edb_top_inst/la0/word_count[9] ), .I2(\edb_top_inst/n2406 ), 
            .O(\edb_top_inst/n2408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3767 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3768  (.I0(\edb_top_inst/edb_user_dr[39] ), 
            .I1(\edb_top_inst/la0/word_count[10] ), .I2(\edb_top_inst/n2408 ), 
            .I3(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3768 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3769  (.I0(\edb_top_inst/la0/word_count[10] ), 
            .I1(\edb_top_inst/n2408 ), .I2(\edb_top_inst/la0/word_count[11] ), 
            .O(\edb_top_inst/n2409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3769 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__3770  (.I0(\edb_top_inst/n2409 ), .I1(\edb_top_inst/edb_user_dr[40] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3770 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3771  (.I0(\edb_top_inst/la0/word_count[10] ), 
            .I1(\edb_top_inst/la0/word_count[11] ), .I2(\edb_top_inst/n2408 ), 
            .O(\edb_top_inst/n2410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3771 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3772  (.I0(\edb_top_inst/edb_user_dr[41] ), 
            .I1(\edb_top_inst/la0/word_count[12] ), .I2(\edb_top_inst/n2410 ), 
            .I3(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3772 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3773  (.I0(\edb_top_inst/la0/word_count[12] ), 
            .I1(\edb_top_inst/n2410 ), .I2(\edb_top_inst/la0/word_count[13] ), 
            .O(\edb_top_inst/n2411 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3773 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__3774  (.I0(\edb_top_inst/n2411 ), .I1(\edb_top_inst/edb_user_dr[42] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3774 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3775  (.I0(\edb_top_inst/la0/word_count[12] ), 
            .I1(\edb_top_inst/la0/word_count[13] ), .I2(\edb_top_inst/n2410 ), 
            .O(\edb_top_inst/n2412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3775 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__3776  (.I0(\edb_top_inst/edb_user_dr[43] ), 
            .I1(\edb_top_inst/la0/word_count[14] ), .I2(\edb_top_inst/n2412 ), 
            .I3(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haa3c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3776 .LUTMASK = 16'haa3c;
    EFX_LUT4 \edb_top_inst/LUT__3777  (.I0(\edb_top_inst/la0/word_count[14] ), 
            .I1(\edb_top_inst/n2412 ), .I2(\edb_top_inst/la0/word_count[15] ), 
            .O(\edb_top_inst/n2413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3777 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__3778  (.I0(\edb_top_inst/n2413 ), .I1(\edb_top_inst/edb_user_dr[44] ), 
            .I2(\edb_top_inst/n2322 ), .O(\edb_top_inst/la0/data_to_word_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3778 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__3779  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n2414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb8f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3779 .LUTMASK = 16'hfb8f;
    EFX_LUT4 \edb_top_inst/LUT__3780  (.I0(\edb_top_inst/n2414 ), .I1(\edb_top_inst/la0/la_trig_mask[1] ), 
            .I2(\edb_top_inst/la0/internal_register_select[3] ), .I3(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n2415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3780 .LUTMASK = 16'h030a;
    EFX_LUT4 \edb_top_inst/LUT__3781  (.I0(\edb_top_inst/n2415 ), .I1(\edb_top_inst/n2367 ), 
            .I2(\edb_top_inst/la0/data_from_biu[1] ), .I3(\edb_top_inst/n2372 ), 
            .O(\edb_top_inst/n2416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3781 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__3782  (.I0(\edb_top_inst/n2416 ), .I1(\edb_top_inst/la0/data_out_shift_reg[2] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3782 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3783  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n2417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3783 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__3784  (.I0(\edb_top_inst/n2417 ), .I1(\edb_top_inst/la0/la_trig_mask[2] ), 
            .I2(\edb_top_inst/la0/internal_register_select[3] ), .I3(\edb_top_inst/la0/internal_register_select[0] ), 
            .O(\edb_top_inst/n2418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3784 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__3785  (.I0(\edb_top_inst/n2418 ), .I1(\edb_top_inst/n2367 ), 
            .I2(\edb_top_inst/la0/data_from_biu[2] ), .I3(\edb_top_inst/n2372 ), 
            .O(\edb_top_inst/n2419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3785 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__3786  (.I0(\edb_top_inst/n2419 ), .I1(\edb_top_inst/la0/data_out_shift_reg[3] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3786 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3787  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/n2372 ), .I2(\edb_top_inst/n2367 ), .O(\edb_top_inst/n2420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3787 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__3788  (.I0(\edb_top_inst/la0/la_sample_cnt[0] ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[3] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3788 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__3789  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[3] ), .I2(\edb_top_inst/n2420 ), 
            .I3(\edb_top_inst/n2421 ), .O(\edb_top_inst/n2422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3789 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__3790  (.I0(\edb_top_inst/n2422 ), .I1(\edb_top_inst/la0/data_out_shift_reg[4] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3790 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3792  (.I0(\edb_top_inst/n2367 ), .I1(\edb_top_inst/la0/internal_register_select[0] ), 
            .I2(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3792 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__3532  (.I0(\edb_top_inst/la0/crc_data_out[6] ), 
            .I1(\edb_top_inst/edb_user_dr[56] ), .I2(\edb_top_inst/la0/crc_data_out[15] ), 
            .I3(\edb_top_inst/edb_user_dr[65] ), .O(\edb_top_inst/n2269 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3532 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3793  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[4] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3793 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__3794  (.I0(\edb_top_inst/n2368 ), .I1(\edb_top_inst/la0/la_trig_mask[4] ), 
            .I2(\edb_top_inst/n2424 ), .I3(\edb_top_inst/n2425 ), .O(\edb_top_inst/n2426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3794 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__3795  (.I0(\edb_top_inst/n2426 ), .I1(\edb_top_inst/la0/data_out_shift_reg[5] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3795 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3796  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[5] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3796 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__3797  (.I0(\edb_top_inst/n2368 ), .I1(\edb_top_inst/la0/la_trig_mask[5] ), 
            .I2(\edb_top_inst/n2424 ), .I3(\edb_top_inst/n2427 ), .O(\edb_top_inst/n2428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3797 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__3798  (.I0(\edb_top_inst/n2428 ), .I1(\edb_top_inst/la0/data_out_shift_reg[6] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3798 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3799  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[6] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3799 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__3800  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[6] ), .I2(\edb_top_inst/n2420 ), 
            .I3(\edb_top_inst/n2429 ), .O(\edb_top_inst/n2430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3800 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__3801  (.I0(\edb_top_inst/n2430 ), .I1(\edb_top_inst/la0/data_out_shift_reg[7] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3801 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3802  (.I0(\edb_top_inst/n2369 ), .I1(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[7] ), .I3(\edb_top_inst/n2368 ), 
            .O(\edb_top_inst/n2431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3802 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3803  (.I0(\edb_top_inst/n2431 ), .I1(\edb_top_inst/la0/data_from_biu[7] ), 
            .I2(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3803 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3804  (.I0(\edb_top_inst/n2432 ), .I1(\edb_top_inst/la0/data_out_shift_reg[8] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3804 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3805  (.I0(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[8] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3805 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__3806  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[8] ), .I2(\edb_top_inst/n2420 ), 
            .I3(\edb_top_inst/n2433 ), .O(\edb_top_inst/n2434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3806 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__3807  (.I0(\edb_top_inst/n2434 ), .I1(\edb_top_inst/la0/data_out_shift_reg[9] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3807 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3808  (.I0(\edb_top_inst/n2369 ), .I1(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[9] ), .I3(\edb_top_inst/n2368 ), 
            .O(\edb_top_inst/n2435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3808 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3809  (.I0(\edb_top_inst/n2435 ), .I1(\edb_top_inst/la0/data_from_biu[9] ), 
            .I2(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3809 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3810  (.I0(\edb_top_inst/n2436 ), .I1(\edb_top_inst/la0/data_out_shift_reg[10] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3810 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3811  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[10] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3811 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__3812  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[10] ), .I2(\edb_top_inst/n2420 ), 
            .I3(\edb_top_inst/n2437 ), .O(\edb_top_inst/n2438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3812 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__3813  (.I0(\edb_top_inst/n2438 ), .I1(\edb_top_inst/la0/data_out_shift_reg[11] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3813 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3814  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[11] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3814 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__3815  (.I0(\edb_top_inst/n2368 ), .I1(\edb_top_inst/la0/la_trig_mask[11] ), 
            .I2(\edb_top_inst/n2424 ), .I3(\edb_top_inst/n2439 ), .O(\edb_top_inst/n2440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3815 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__3816  (.I0(\edb_top_inst/n2440 ), .I1(\edb_top_inst/la0/data_out_shift_reg[12] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3816 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3817  (.I0(\edb_top_inst/n2369 ), .I1(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[12] ), .I3(\edb_top_inst/n2368 ), 
            .O(\edb_top_inst/n2441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3817 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3818  (.I0(\edb_top_inst/n2441 ), .I1(\edb_top_inst/la0/data_from_biu[12] ), 
            .I2(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3818 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3819  (.I0(\edb_top_inst/n2442 ), .I1(\edb_top_inst/la0/data_out_shift_reg[13] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3819 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3820  (.I0(\edb_top_inst/n2369 ), .I1(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[13] ), .I3(\edb_top_inst/n2368 ), 
            .O(\edb_top_inst/n2443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3820 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3821  (.I0(\edb_top_inst/n2443 ), .I1(\edb_top_inst/la0/data_from_biu[13] ), 
            .I2(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3821 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3822  (.I0(\edb_top_inst/n2444 ), .I1(\edb_top_inst/la0/data_out_shift_reg[14] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3822 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3823  (.I0(\edb_top_inst/la0/la_sample_cnt[11] ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[14] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3823 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__3824  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[14] ), .I2(\edb_top_inst/n2420 ), 
            .I3(\edb_top_inst/n2445 ), .O(\edb_top_inst/n2446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3824 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__3825  (.I0(\edb_top_inst/n2446 ), .I1(\edb_top_inst/la0/data_out_shift_reg[15] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3825 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3826  (.I0(\edb_top_inst/la0/la_trig_mask[15] ), 
            .I1(\edb_top_inst/n2368 ), .I2(\edb_top_inst/la0/data_from_biu[15] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3826 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__3827  (.I0(\edb_top_inst/n2447 ), .I1(\edb_top_inst/la0/data_out_shift_reg[16] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3827 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3828  (.I0(\edb_top_inst/la0/la_trig_mask[16] ), 
            .I1(\edb_top_inst/n2368 ), .I2(\edb_top_inst/la0/data_from_biu[16] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3828 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__3829  (.I0(\edb_top_inst/n2448 ), .I1(\edb_top_inst/la0/data_out_shift_reg[17] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3829 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3830  (.I0(\edb_top_inst/la0/la_trig_mask[17] ), 
            .I1(\edb_top_inst/la0/internal_register_select[0] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/n2367 ), .O(\edb_top_inst/n2449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3830 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__3831  (.I0(\edb_top_inst/n2449 ), .I1(\edb_top_inst/la0/data_from_biu[17] ), 
            .I2(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3831 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3832  (.I0(\edb_top_inst/n2450 ), .I1(\edb_top_inst/la0/data_out_shift_reg[18] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3832 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3833  (.I0(\edb_top_inst/la0/la_trig_mask[18] ), 
            .I1(\edb_top_inst/n2368 ), .I2(\edb_top_inst/la0/data_from_biu[18] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3833 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__3834  (.I0(\edb_top_inst/n2451 ), .I1(\edb_top_inst/la0/data_out_shift_reg[19] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3834 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3835  (.I0(\edb_top_inst/la0/la_trig_mask[19] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/la0/internal_register_select[0] ), 
            .I3(\edb_top_inst/n2367 ), .O(\edb_top_inst/n2452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3835 .LUTMASK = 16'h2c00;
    EFX_LUT4 \edb_top_inst/LUT__3836  (.I0(\edb_top_inst/n2452 ), .I1(\edb_top_inst/la0/data_from_biu[19] ), 
            .I2(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3836 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3837  (.I0(\edb_top_inst/n2453 ), .I1(\edb_top_inst/la0/data_out_shift_reg[20] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3837 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3838  (.I0(\edb_top_inst/la0/la_run_trig ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[20] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3838 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__3839  (.I0(\edb_top_inst/n2368 ), .I1(\edb_top_inst/la0/la_trig_mask[20] ), 
            .I2(\edb_top_inst/n2424 ), .I3(\edb_top_inst/n2454 ), .O(\edb_top_inst/n2455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3839 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__3840  (.I0(\edb_top_inst/n2455 ), .I1(\edb_top_inst/la0/data_out_shift_reg[21] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3840 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3841  (.I0(\edb_top_inst/la0/la_run_trig_imdt ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[21] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3841 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__3842  (.I0(\edb_top_inst/n2368 ), .I1(\edb_top_inst/la0/la_trig_mask[21] ), 
            .I2(\edb_top_inst/n2424 ), .I3(\edb_top_inst/n2456 ), .O(\edb_top_inst/n2457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3842 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__3843  (.I0(\edb_top_inst/n2457 ), .I1(\edb_top_inst/la0/data_out_shift_reg[22] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3843 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3844  (.I0(\edb_top_inst/la0/la_stop_trig ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[22] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3844 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__3845  (.I0(\edb_top_inst/n2368 ), .I1(\edb_top_inst/la0/la_trig_mask[22] ), 
            .I2(\edb_top_inst/n2424 ), .I3(\edb_top_inst/n2458 ), .O(\edb_top_inst/n2459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3845 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__3846  (.I0(\edb_top_inst/n2459 ), .I1(\edb_top_inst/la0/data_out_shift_reg[23] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3846 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3847  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[23] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3847 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__3848  (.I0(\edb_top_inst/n2368 ), .I1(\edb_top_inst/la0/la_trig_mask[23] ), 
            .I2(\edb_top_inst/n2424 ), .I3(\edb_top_inst/n2460 ), .O(\edb_top_inst/n2461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3848 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__3849  (.I0(\edb_top_inst/n2461 ), .I1(\edb_top_inst/la0/data_out_shift_reg[24] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3849 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3850  (.I0(\edb_top_inst/n2369 ), .I1(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[24] ), .I3(\edb_top_inst/n2368 ), 
            .O(\edb_top_inst/n2462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3850 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3851  (.I0(\edb_top_inst/n2462 ), .I1(\edb_top_inst/la0/data_from_biu[24] ), 
            .I2(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2463 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3851 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3852  (.I0(\edb_top_inst/n2463 ), .I1(\edb_top_inst/la0/data_out_shift_reg[25] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3852 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3853  (.I0(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[25] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3853 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__3854  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[25] ), .I2(\edb_top_inst/n2420 ), 
            .I3(\edb_top_inst/n2464 ), .O(\edb_top_inst/n2465 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3854 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__3855  (.I0(\edb_top_inst/n2465 ), .I1(\edb_top_inst/la0/data_out_shift_reg[26] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3855 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3856  (.I0(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[26] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3856 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__3857  (.I0(\edb_top_inst/n2466 ), .I1(\edb_top_inst/n2367 ), 
            .I2(\edb_top_inst/la0/data_from_biu[26] ), .I3(\edb_top_inst/n2372 ), 
            .O(\edb_top_inst/n2467 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3857 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__3858  (.I0(\edb_top_inst/n2467 ), .I1(\edb_top_inst/la0/data_out_shift_reg[27] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3858 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3859  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[27] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3859 .LUTMASK = 16'hbbf0;
    EFX_LUT4 \edb_top_inst/LUT__3860  (.I0(\edb_top_inst/n2368 ), .I1(\edb_top_inst/la0/la_trig_mask[27] ), 
            .I2(\edb_top_inst/n2424 ), .I3(\edb_top_inst/n2468 ), .O(\edb_top_inst/n2469 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3860 .LUTMASK = 16'h8f00;
    EFX_LUT4 \edb_top_inst/LUT__3861  (.I0(\edb_top_inst/n2469 ), .I1(\edb_top_inst/la0/data_out_shift_reg[28] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3861 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3862  (.I0(\edb_top_inst/n2369 ), .I1(\edb_top_inst/la0/la_trig_pos[5] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[28] ), .I3(\edb_top_inst/n2368 ), 
            .O(\edb_top_inst/n2470 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3862 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3863  (.I0(\edb_top_inst/n2470 ), .I1(\edb_top_inst/la0/data_from_biu[28] ), 
            .I2(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2471 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3863 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3864  (.I0(\edb_top_inst/n2471 ), .I1(\edb_top_inst/la0/data_out_shift_reg[29] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3864 .LUTMASK = 16'hacac;
    EFX_LUT4 \edb_top_inst/LUT__3865  (.I0(\edb_top_inst/la0/la_trig_pos[6] ), 
            .I1(\edb_top_inst/n2369 ), .I2(\edb_top_inst/la0/data_from_biu[29] ), 
            .I3(\edb_top_inst/n2372 ), .O(\edb_top_inst/n2472 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3865 .LUTMASK = 16'h770f;
    EFX_LUT4 \edb_top_inst/LUT__3866  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[29] ), .I2(\edb_top_inst/n2420 ), 
            .I3(\edb_top_inst/n2472 ), .O(\edb_top_inst/n2473 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3866 .LUTMASK = 16'h1f00;
    EFX_LUT4 \edb_top_inst/LUT__3867  (.I0(\edb_top_inst/n2473 ), .I1(\edb_top_inst/la0/data_out_shift_reg[30] ), 
            .I2(\edb_top_inst/n2375 ), .O(\edb_top_inst/la0/n2431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c5c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3867 .LUTMASK = 16'h5c5c;
    EFX_LUT4 \edb_top_inst/LUT__3868  (.I0(\edb_top_inst/n2369 ), .I1(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[30] ), .I3(\edb_top_inst/n2368 ), 
            .O(\edb_top_inst/n2474 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3868 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3869  (.I0(\edb_top_inst/n2474 ), .I1(\edb_top_inst/n2372 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[31] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3869 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3870  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[31] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2475 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3870 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__3871  (.I0(\edb_top_inst/n2372 ), .I1(\edb_top_inst/n2367 ), 
            .O(\edb_top_inst/n2476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3871 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__3872  (.I0(\edb_top_inst/n2476 ), .I1(\edb_top_inst/n2475 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[32] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3872 .LUTMASK = 16'h88f0;
    EFX_LUT4 \edb_top_inst/LUT__3873  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[32] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2477 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3873 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__3874  (.I0(\edb_top_inst/n2476 ), .I1(\edb_top_inst/n2477 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[33] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3874 .LUTMASK = 16'h88f0;
    EFX_LUT4 \edb_top_inst/LUT__3875  (.I0(\edb_top_inst/n2369 ), .I1(\edb_top_inst/la0/la_trig_pos[10] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[33] ), .I3(\edb_top_inst/n2368 ), 
            .O(\edb_top_inst/n2478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3875 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3876  (.I0(\edb_top_inst/n2478 ), .I1(\edb_top_inst/n2372 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[34] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3876 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3877  (.I0(\edb_top_inst/la0/la_trig_mask[34] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[11] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2479 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3877 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__3878  (.I0(\edb_top_inst/n2476 ), .I1(\edb_top_inst/n2479 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[35] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3878 .LUTMASK = 16'h88f0;
    EFX_LUT4 \edb_top_inst/LUT__3879  (.I0(\edb_top_inst/la0/la_trig_pos[12] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[35] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3879 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__3880  (.I0(\edb_top_inst/n2476 ), .I1(\edb_top_inst/n2480 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[36] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3880 .LUTMASK = 16'h88f0;
    EFX_LUT4 \edb_top_inst/LUT__3881  (.I0(\edb_top_inst/la0/la_trig_pos[13] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[36] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2481 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3881 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__3882  (.I0(\edb_top_inst/n2481 ), .I1(\edb_top_inst/n2476 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[37] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3882 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3883  (.I0(\edb_top_inst/la0/la_trig_pos[14] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[37] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2482 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3883 .LUTMASK = 16'h0305;
    EFX_LUT4 \edb_top_inst/LUT__3884  (.I0(\edb_top_inst/n2482 ), .I1(\edb_top_inst/n2476 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[38] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2423 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3884 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3885  (.I0(\edb_top_inst/n2369 ), .I1(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[38] ), .I3(\edb_top_inst/n2368 ), 
            .O(\edb_top_inst/n2483 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3885 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3886  (.I0(\edb_top_inst/n2483 ), .I1(\edb_top_inst/n2372 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[39] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3886 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3887  (.I0(\edb_top_inst/la0/la_trig_mask[39] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[16] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2484 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0afc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3887 .LUTMASK = 16'h0afc;
    EFX_LUT4 \edb_top_inst/LUT__3888  (.I0(\edb_top_inst/n2476 ), .I1(\edb_top_inst/n2484 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[40] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3888 .LUTMASK = 16'h88f0;
    EFX_LUT4 \edb_top_inst/LUT__3889  (.I0(\edb_top_inst/la0/la_trig_mask[40] ), 
            .I1(\edb_top_inst/n2368 ), .I2(\edb_top_inst/la0/la_trig_pattern[0] ), 
            .I3(\edb_top_inst/n2369 ), .O(\edb_top_inst/n2485 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3889 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3890  (.I0(\edb_top_inst/n2485 ), .I1(\edb_top_inst/n2372 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[41] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3890 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3891  (.I0(\edb_top_inst/la0/la_trig_pattern[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[41] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2486 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3891 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__3892  (.I0(\edb_top_inst/n2476 ), .I1(\edb_top_inst/n2486 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[42] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3892 .LUTMASK = 16'h88f0;
    EFX_LUT4 \edb_top_inst/LUT__3893  (.I0(\edb_top_inst/la0/la_trig_mask[42] ), 
            .I1(\edb_top_inst/n2368 ), .I2(\edb_top_inst/la0/la_capture_pattern[0] ), 
            .I3(\edb_top_inst/n2369 ), .O(\edb_top_inst/n2487 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3893 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__3894  (.I0(\edb_top_inst/n2487 ), .I1(\edb_top_inst/n2372 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[43] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3894 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3895  (.I0(\edb_top_inst/la0/la_capture_pattern[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[43] ), .I2(\edb_top_inst/la0/internal_register_select[3] ), 
            .I3(\edb_top_inst/la0/internal_register_select[0] ), .O(\edb_top_inst/n2488 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3895 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__3896  (.I0(\edb_top_inst/n2476 ), .I1(\edb_top_inst/n2488 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[44] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3896 .LUTMASK = 16'h88f0;
    EFX_LUT4 \edb_top_inst/LUT__3897  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/n2372 ), 
            .I2(\edb_top_inst/n2368 ), .O(\edb_top_inst/n2489 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3897 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__3898  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/la0/data_out_shift_reg[45] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[44] ), .I3(\edb_top_inst/n2489 ), 
            .O(\edb_top_inst/la0/n2416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3898 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3899  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/la0/data_out_shift_reg[46] ), 
            .O(\edb_top_inst/n2490 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3899 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3900  (.I0(\edb_top_inst/la0/internal_register_select[0] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .I2(\edb_top_inst/n2375 ), 
            .I3(\edb_top_inst/n2476 ), .O(\edb_top_inst/n2491 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3900 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__3901  (.I0(\edb_top_inst/n2489 ), .I1(\edb_top_inst/la0/la_trig_mask[45] ), 
            .I2(\edb_top_inst/n2490 ), .I3(\edb_top_inst/n2491 ), .O(\edb_top_inst/la0/n2415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3901 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__3902  (.I0(\edb_top_inst/la0/la_trig_mask[46] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n2492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3902 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3903  (.I0(\edb_top_inst/la0/internal_register_select[3] ), 
            .I1(\edb_top_inst/la0/internal_register_select[0] ), .I2(\edb_top_inst/n2375 ), 
            .I3(\edb_top_inst/n2476 ), .O(\edb_top_inst/n2493 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3903 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__3904  (.I0(\edb_top_inst/n2492 ), .I1(\edb_top_inst/n2493 ), 
            .I2(\edb_top_inst/n2375 ), .I3(\edb_top_inst/la0/data_out_shift_reg[47] ), 
            .O(\edb_top_inst/la0/n2414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3904 .LUTMASK = 16'h4f44;
    EFX_LUT4 \edb_top_inst/LUT__3905  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/la0/data_out_shift_reg[48] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[47] ), .I3(\edb_top_inst/n2489 ), 
            .O(\edb_top_inst/la0/n2413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3905 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3906  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/la0/data_out_shift_reg[49] ), 
            .O(\edb_top_inst/n2494 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3906 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3907  (.I0(\edb_top_inst/n2489 ), .I1(\edb_top_inst/la0/la_trig_mask[48] ), 
            .I2(\edb_top_inst/n2491 ), .I3(\edb_top_inst/n2494 ), .O(\edb_top_inst/la0/n2412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3907 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__3908  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/la0/data_out_shift_reg[50] ), 
            .O(\edb_top_inst/n2495 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3908 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3909  (.I0(\edb_top_inst/n2489 ), .I1(\edb_top_inst/la0/la_trig_mask[49] ), 
            .I2(\edb_top_inst/n2491 ), .I3(\edb_top_inst/n2495 ), .O(\edb_top_inst/la0/n2411 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3909 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__3910  (.I0(\edb_top_inst/la0/la_trig_mask[50] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n2496 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3910 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3911  (.I0(\edb_top_inst/n2496 ), .I1(\edb_top_inst/n2493 ), 
            .I2(\edb_top_inst/n2375 ), .I3(\edb_top_inst/la0/data_out_shift_reg[51] ), 
            .O(\edb_top_inst/la0/n2410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3911 .LUTMASK = 16'h4f44;
    EFX_LUT4 \edb_top_inst/LUT__3912  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/la0/data_out_shift_reg[52] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[51] ), .I3(\edb_top_inst/n2489 ), 
            .O(\edb_top_inst/la0/n2409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3912 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3913  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/la0/data_out_shift_reg[53] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[52] ), .I3(\edb_top_inst/n2489 ), 
            .O(\edb_top_inst/la0/n2408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3913 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3914  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/la0/data_out_shift_reg[54] ), 
            .O(\edb_top_inst/n2497 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3914 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3915  (.I0(\edb_top_inst/n2489 ), .I1(\edb_top_inst/la0/la_trig_mask[53] ), 
            .I2(\edb_top_inst/n2491 ), .I3(\edb_top_inst/n2497 ), .O(\edb_top_inst/la0/n2407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3915 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__3916  (.I0(\edb_top_inst/la0/la_trig_mask[54] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n2498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3916 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3917  (.I0(\edb_top_inst/n2498 ), .I1(\edb_top_inst/n2420 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[55] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3917 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3918  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/la0/data_out_shift_reg[56] ), 
            .O(\edb_top_inst/n2499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3918 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3919  (.I0(\edb_top_inst/n2489 ), .I1(\edb_top_inst/la0/la_trig_mask[55] ), 
            .I2(\edb_top_inst/n2491 ), .I3(\edb_top_inst/n2499 ), .O(\edb_top_inst/la0/n2405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3919 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__3920  (.I0(\edb_top_inst/la0/la_trig_mask[56] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n2500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3920 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3921  (.I0(\edb_top_inst/n2500 ), .I1(\edb_top_inst/n2420 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[57] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3921 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3922  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/la0/data_out_shift_reg[58] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[57] ), .I3(\edb_top_inst/n2489 ), 
            .O(\edb_top_inst/la0/n2403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3922 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3923  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/la0/data_out_shift_reg[59] ), 
            .O(\edb_top_inst/n2501 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3923 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__3924  (.I0(\edb_top_inst/n2489 ), .I1(\edb_top_inst/la0/la_trig_mask[58] ), 
            .I2(\edb_top_inst/n2491 ), .I3(\edb_top_inst/n2501 ), .O(\edb_top_inst/la0/n2402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3924 .LUTMASK = 16'hfff8;
    EFX_LUT4 \edb_top_inst/LUT__3925  (.I0(\edb_top_inst/la0/la_trig_mask[59] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n2502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3925 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3926  (.I0(\edb_top_inst/n2502 ), .I1(\edb_top_inst/n2493 ), 
            .I2(\edb_top_inst/n2375 ), .I3(\edb_top_inst/la0/data_out_shift_reg[60] ), 
            .O(\edb_top_inst/la0/n2401 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3926 .LUTMASK = 16'h4f44;
    EFX_LUT4 \edb_top_inst/LUT__3927  (.I0(\edb_top_inst/la0/la_trig_mask[60] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n2503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3927 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3928  (.I0(\edb_top_inst/n2503 ), .I1(\edb_top_inst/n2420 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[61] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2400 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3928 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3929  (.I0(\edb_top_inst/n2375 ), .I1(\edb_top_inst/la0/data_out_shift_reg[62] ), 
            .I2(\edb_top_inst/la0/la_trig_mask[61] ), .I3(\edb_top_inst/n2489 ), 
            .O(\edb_top_inst/la0/n2399 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3929 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__3930  (.I0(\edb_top_inst/la0/la_trig_mask[62] ), 
            .I1(\edb_top_inst/la0/internal_register_select[3] ), .O(\edb_top_inst/n2504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3930 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__3931  (.I0(\edb_top_inst/n2504 ), .I1(\edb_top_inst/n2420 ), 
            .I2(\edb_top_inst/la0/data_out_shift_reg[63] ), .I3(\edb_top_inst/n2375 ), 
            .O(\edb_top_inst/la0/n2398 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h44f0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3931 .LUTMASK = 16'h44f0;
    EFX_LUT4 \edb_top_inst/LUT__3932  (.I0(\edb_top_inst/n2489 ), .I1(\edb_top_inst/la0/la_trig_mask[63] ), 
            .I2(\edb_top_inst/n2491 ), .O(\edb_top_inst/la0/n2397 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3932 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__3933  (.I0(\edb_top_inst/n2344 ), .I1(\edb_top_inst/n2358 ), 
            .I2(jtag_inst1_UPDATE), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n2505 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3933 .LUTMASK = 16'h7077;
    EFX_LUT4 \edb_top_inst/LUT__3934  (.I0(\edb_top_inst/n2312 ), .I1(\edb_top_inst/n2343 ), 
            .I2(\edb_top_inst/la0/module_state[0] ), .I3(\edb_top_inst/la0/module_state[1] ), 
            .O(\edb_top_inst/n2506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf50, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3934 .LUTMASK = 16'hcf50;
    EFX_LUT4 \edb_top_inst/LUT__3935  (.I0(\edb_top_inst/n2506 ), .I1(\edb_top_inst/n2505 ), 
            .I2(\edb_top_inst/la0/module_state[3] ), .I3(\edb_top_inst/la0/module_state[2] ), 
            .O(\edb_top_inst/n2507 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3935 .LUTMASK = 16'h030a;
    EFX_LUT4 \edb_top_inst/LUT__3936  (.I0(\edb_top_inst/n2357 ), .I1(jtag_inst1_UPDATE), 
            .I2(\edb_top_inst/n2293 ), .I3(\edb_top_inst/n2507 ), .O(\edb_top_inst/la0/module_next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3936 .LUTMASK = 16'hff10;
    EFX_LUT4 \edb_top_inst/LUT__3937  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/n2304 ), .I2(\edb_top_inst/n2355 ), .I3(\edb_top_inst/n2312 ), 
            .O(\edb_top_inst/n2508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3937 .LUTMASK = 16'he800;
    EFX_LUT4 \edb_top_inst/LUT__3938  (.I0(\edb_top_inst/n2357 ), .I1(jtag_inst1_UPDATE), 
            .I2(\edb_top_inst/n2305 ), .O(\edb_top_inst/n2509 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3938 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__3939  (.I0(jtag_inst1_UPDATE), .I1(\edb_top_inst/n2312 ), 
            .I2(\edb_top_inst/n2293 ), .I3(\edb_top_inst/n2307 ), .O(\edb_top_inst/n2510 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3939 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__3940  (.I0(\edb_top_inst/n2509 ), .I1(\edb_top_inst/n2508 ), 
            .I2(\edb_top_inst/n2356 ), .I3(\edb_top_inst/n2510 ), .O(\edb_top_inst/la0/module_next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3940 .LUTMASK = 16'hfff2;
    EFX_LUT4 \edb_top_inst/LUT__3941  (.I0(\edb_top_inst/la0/crc_data_out[1] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3941 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3942  (.I0(\edb_top_inst/n2357 ), .I1(\edb_top_inst/n2293 ), 
            .I2(\edb_top_inst/la0/op_reg_en ), .I3(\edb_top_inst/n2363 ), 
            .O(\edb_top_inst/ceg_net221 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3942 .LUTMASK = 16'h0007;
    EFX_LUT4 \edb_top_inst/LUT__3943  (.I0(\edb_top_inst/la0/crc_data_out[2] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n149 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3943 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3944  (.I0(\edb_top_inst/la0/crc_data_out[3] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3944 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3945  (.I0(\edb_top_inst/la0/crc_data_out[4] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n147 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3945 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3946  (.I0(\edb_top_inst/la0/crc_data_out[5] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3946 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3947  (.I0(jtag_inst1_TDI), .I1(\edb_top_inst/la0/data_out_shift_reg[0] ), 
            .I2(\edb_top_inst/la0/module_state[1] ), .I3(\edb_top_inst/la0/crc_data_out[0] ), 
            .O(\edb_top_inst/n2511 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h53ac, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3947 .LUTMASK = 16'h53ac;
    EFX_LUT4 \edb_top_inst/LUT__3948  (.I0(\edb_top_inst/n2357 ), .I1(\edb_top_inst/n2511 ), 
            .I2(\edb_top_inst/n2305 ), .O(\edb_top_inst/n2512 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3948 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__3949  (.I0(\edb_top_inst/la0/module_state[0] ), 
            .I1(\edb_top_inst/n2350 ), .I2(\edb_top_inst/la0/module_state[1] ), 
            .I3(\edb_top_inst/n2512 ), .O(\edb_top_inst/n2513 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3949 .LUTMASK = 16'hbf00;
    EFX_LUT4 \edb_top_inst/LUT__3950  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[6] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n145 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3950 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3951  (.I0(\edb_top_inst/la0/crc_data_out[7] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3951 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3952  (.I0(\edb_top_inst/la0/crc_data_out[8] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n143 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3952 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3953  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[9] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3953 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3954  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[10] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n141 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3954 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3955  (.I0(\edb_top_inst/la0/crc_data_out[11] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3955 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3956  (.I0(\edb_top_inst/la0/crc_data_out[12] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n139 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3956 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3957  (.I0(\edb_top_inst/la0/crc_data_out[13] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3957 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3958  (.I0(\edb_top_inst/la0/crc_data_out[14] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3958 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3959  (.I0(\edb_top_inst/la0/crc_data_out[15] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3959 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3960  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[16] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n135 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3960 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3961  (.I0(\edb_top_inst/la0/crc_data_out[17] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3961 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3962  (.I0(\edb_top_inst/la0/crc_data_out[18] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n133 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3962 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3963  (.I0(\edb_top_inst/la0/crc_data_out[19] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3963 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3964  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[20] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n131 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3964 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3965  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[21] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3965 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3966  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[22] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n129 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3966 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3967  (.I0(\edb_top_inst/la0/crc_data_out[23] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3967 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3968  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[24] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n127 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3968 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3969  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[25] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3969 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3970  (.I0(\edb_top_inst/la0/crc_data_out[26] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n125 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3970 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3971  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[27] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3971 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3972  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[28] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n123 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3972 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3973  (.I0(\edb_top_inst/la0/crc_data_out[29] ), 
            .I1(\edb_top_inst/la0/op_reg_en ), .O(\edb_top_inst/la0/axi_crc_i/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3973 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3974  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[30] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3974 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3975  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/la0/crc_data_out[31] ), .I2(\edb_top_inst/n2513 ), 
            .O(\edb_top_inst/la0/axi_crc_i/n120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3975 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__3976  (.I0(\edb_top_inst/la0/op_reg_en ), 
            .I1(\edb_top_inst/n2513 ), .O(\edb_top_inst/la0/axi_crc_i/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3976 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__3977  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3977 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3978  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3978 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3979  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b22, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3979 .LUTMASK = 16'h2b22;
    EFX_LUT4 \edb_top_inst/LUT__3980  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/equal_9/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ff6, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3980 .LUTMASK = 16'h6ff6;
    EFX_LUT4 \edb_top_inst/LUT__3981  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n2514 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3981 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__3982  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/n2514 ), .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n2515 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3982 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__3983  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n2516 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3983 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3984  (.I0(\edb_top_inst/n2514 ), .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n2516 ), .O(\edb_top_inst/n2517 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4c70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3984 .LUTMASK = 16'h4c70;
    EFX_LUT4 \edb_top_inst/LUT__3985  (.I0(\edb_top_inst/n2517 ), .I1(\edb_top_inst/n2515 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3985 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__3986  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3986 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3987  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.capture_cu/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3987 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3988  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3988 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3989  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3989 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3990  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b22, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3990 .LUTMASK = 16'h2b22;
    EFX_LUT4 \edb_top_inst/LUT__3991  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/equal_9/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ff6, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3991 .LUTMASK = 16'h6ff6;
    EFX_LUT4 \edb_top_inst/LUT__3992  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n2518 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3992 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__3993  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/n2518 ), .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n2519 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3993 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__3994  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n2520 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3994 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__3995  (.I0(\edb_top_inst/n2518 ), .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n2520 ), .O(\edb_top_inst/n2521 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4c70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3995 .LUTMASK = 16'h4c70;
    EFX_LUT4 \edb_top_inst/LUT__3996  (.I0(\edb_top_inst/n2521 ), .I1(\edb_top_inst/n2519 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3996 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__3997  (.I0(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3997 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3998  (.I0(\edb_top_inst/la0/GEN_PROBE[0].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[0].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.trigger_cu/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3998 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__3999  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n2522 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__3999 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__4000  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n2522 ), .O(\edb_top_inst/n2523 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4000 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__4001  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n2524 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4001 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4002  (.I0(\edb_top_inst/n2524 ), .I1(\edb_top_inst/n2523 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4002 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4003  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/genblk1.rise )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4003 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4004  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/genblk1.fall )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4004 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4005  (.I0(\edb_top_inst/la0/GEN_PROBE[1].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4005 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4006  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/n18 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.enable ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.capture_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4006 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4007  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp6 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp5 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n2525 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha0cf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4007 .LUTMASK = 16'ha0cf;
    EFX_LUT4 \edb_top_inst/LUT__4008  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp4 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp3 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n2525 ), .O(\edb_top_inst/n2526 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfc0a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4008 .LUTMASK = 16'hfc0a;
    EFX_LUT4 \edb_top_inst/LUT__4009  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.data_in_p1 ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n2527 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4009 .LUTMASK = 16'hfac0;
    EFX_LUT4 \edb_top_inst/LUT__4010  (.I0(\edb_top_inst/n2527 ), .I1(\edb_top_inst/n2526 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4010 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4011  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4011 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4012  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4012 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4013  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b22, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4013 .LUTMASK = 16'h2b22;
    EFX_LUT4 \edb_top_inst/LUT__4014  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/equal_9/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ff6, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4014 .LUTMASK = 16'h6ff6;
    EFX_LUT4 \edb_top_inst/LUT__4015  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n2528 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4015 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__4016  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/n2528 ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n2529 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4016 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__4017  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n2530 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4017 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4018  (.I0(\edb_top_inst/n2528 ), .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n2530 ), .O(\edb_top_inst/n2531 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4c70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4018 .LUTMASK = 16'h4c70;
    EFX_LUT4 \edb_top_inst/LUT__4019  (.I0(\edb_top_inst/n2531 ), .I1(\edb_top_inst/n2529 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4019 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4020  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4020 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4021  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.capture_cu/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4021 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4022  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4022 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4023  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n10 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4023 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4024  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b22, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4024 .LUTMASK = 16'h2b22;
    EFX_LUT4 \edb_top_inst/LUT__4025  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/equal_9/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6ff6, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4025 .LUTMASK = 16'h6ff6;
    EFX_LUT4 \edb_top_inst/LUT__4026  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n2532 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4026 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__4027  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/n2532 ), .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/n2533 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4027 .LUTMASK = 16'he3e3;
    EFX_LUT4 \edb_top_inst/LUT__4028  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n2534 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4028 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4029  (.I0(\edb_top_inst/n2532 ), .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/n2534 ), .O(\edb_top_inst/n2535 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h704c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4029 .LUTMASK = 16'h704c;
    EFX_LUT4 \edb_top_inst/LUT__4030  (.I0(\edb_top_inst/n2535 ), .I1(\edb_top_inst/n2533 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4030 .LUTMASK = 16'h3a3a;
    EFX_LUT4 \edb_top_inst/LUT__4031  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4031 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4032  (.I0(\edb_top_inst/la0/GEN_PROBE[2].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.trigger_cu/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4032 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4033  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4033 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4034  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4034 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4035  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), .O(\edb_top_inst/n2536 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4035 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4036  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/n2536 ), .O(\edb_top_inst/n2537 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4036 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__4037  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/n2537 ), .O(\edb_top_inst/n2538 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4037 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4038  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/n2538 ), .O(\edb_top_inst/n2539 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4038 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4039  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/n2539 ), .O(\edb_top_inst/n2540 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4039 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4040  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/n2541 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4040 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4041  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9] ), .O(\edb_top_inst/n2542 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4041 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4042  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11] ), .O(\edb_top_inst/n2543 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4042 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4043  (.I0(\edb_top_inst/n2542 ), .I1(\edb_top_inst/n2541 ), 
            .I2(\edb_top_inst/n2543 ), .O(\edb_top_inst/n2544 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4043 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4044  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7] ), .O(\edb_top_inst/n2545 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4044 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4045  (.I0(\edb_top_inst/n2544 ), .I1(\edb_top_inst/n2545 ), 
            .O(\edb_top_inst/n2546 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4045 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4046  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6] ), 
            .I1(\edb_top_inst/n2540 ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/n2546 ), .O(\edb_top_inst/n2547 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4046 .LUTMASK = 16'h7100;
    EFX_LUT4 \edb_top_inst/LUT__4047  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n2548 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4047 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__4048  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/n2549 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4048 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4049  (.I0(\edb_top_inst/n2548 ), .I1(\edb_top_inst/n2541 ), 
            .I2(\edb_top_inst/n2549 ), .I3(\edb_top_inst/n2544 ), .O(\edb_top_inst/n2550 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4049 .LUTMASK = 16'hbf00;
    EFX_LUT4 \edb_top_inst/LUT__4050  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/n2551 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4050 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4051  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n2552 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4051 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4052  (.I0(\edb_top_inst/n2551 ), .I1(\edb_top_inst/n2552 ), 
            .O(\edb_top_inst/n2553 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4052 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4053  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13] ), .O(\edb_top_inst/n2554 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4053 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4054  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15] ), 
            .I2(\edb_top_inst/n2554 ), .O(\edb_top_inst/n2555 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4054 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__4055  (.I0(\edb_top_inst/n2550 ), .I1(\edb_top_inst/n2547 ), 
            .I2(\edb_top_inst/n2553 ), .I3(\edb_top_inst/n2555 ), .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4055 .LUTMASK = 16'hff10;
    EFX_LUT4 \edb_top_inst/LUT__4056  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n2556 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4056 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4057  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n2557 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4057 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4058  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n2558 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4058 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4059  (.I0(\edb_top_inst/n2556 ), .I1(\edb_top_inst/n2552 ), 
            .I2(\edb_top_inst/n2557 ), .I3(\edb_top_inst/n2558 ), .O(\edb_top_inst/n2559 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4059 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4060  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n2560 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4060 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4061  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/n2561 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4061 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4062  (.I0(\edb_top_inst/n2560 ), .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] ), .I3(\edb_top_inst/n2561 ), 
            .O(\edb_top_inst/n2562 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4062 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__4063  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n2563 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4063 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4064  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n2564 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4064 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4065  (.I0(\edb_top_inst/n2559 ), .I1(\edb_top_inst/n2562 ), 
            .I2(\edb_top_inst/n2563 ), .I3(\edb_top_inst/n2564 ), .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/equal_9/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4065 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4066  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n2565 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4066 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4067  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[13] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n2566 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4067 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4068  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[11] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[12] ), 
            .O(\edb_top_inst/n2567 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4068 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4069  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[9] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[10] ), 
            .O(\edb_top_inst/n2568 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4069 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4070  (.I0(\edb_top_inst/n2565 ), .I1(\edb_top_inst/n2566 ), 
            .I2(\edb_top_inst/n2567 ), .I3(\edb_top_inst/n2568 ), .O(\edb_top_inst/n2569 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4070 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4071  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4] ), 
            .O(\edb_top_inst/n2570 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4071 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4072  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n2571 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4072 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4073  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2] ), 
            .O(\edb_top_inst/n2572 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4073 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4074  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6] ), 
            .O(\edb_top_inst/n2573 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4074 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4075  (.I0(\edb_top_inst/n2570 ), .I1(\edb_top_inst/n2571 ), 
            .I2(\edb_top_inst/n2572 ), .I3(\edb_top_inst/n2573 ), .O(\edb_top_inst/n2574 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4075 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4076  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/n2569 ), .I3(\edb_top_inst/n2574 ), .O(\edb_top_inst/n2575 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4076 .LUTMASK = 16'haccc;
    EFX_LUT4 \edb_top_inst/LUT__4077  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n2576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4077 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4078  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n2577 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4078 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__4079  (.I0(\edb_top_inst/n2576 ), .I1(\edb_top_inst/n2575 ), 
            .I2(\edb_top_inst/n2577 ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f44, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4079 .LUTMASK = 16'h0f44;
    EFX_LUT4 \edb_top_inst/LUT__4080  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4080 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4081  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4081 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4082  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4082 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4083  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4083 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4084  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4084 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4085  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4085 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4086  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4086 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4087  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4087 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4088  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4088 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4089  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4089 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4090  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4090 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4091  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4091 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4092  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4092 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4093  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4093 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4094  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4094 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4095  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4095 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4096  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4096 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4097  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4097 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4098  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4098 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4099  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4099 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4100  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4100 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4101  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4101 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4102  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4102 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4103  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4103 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4104  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4104 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4105  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4105 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4106  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4106 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4107  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4107 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4108  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4108 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4109  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.capture_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4109 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4110  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4110 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4111  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4111 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4112  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), .O(\edb_top_inst/n2578 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4112 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4113  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/n2578 ), .O(\edb_top_inst/n2579 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4113 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__4114  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I2(\edb_top_inst/n2579 ), .O(\edb_top_inst/n2580 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4114 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4115  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/n2580 ), .O(\edb_top_inst/n2581 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4115 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4116  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/n2581 ), .O(\edb_top_inst/n2582 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4116 .LUTMASK = 16'hb2b2;
    EFX_LUT4 \edb_top_inst/LUT__4117  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/n2583 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4117 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4118  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9] ), .O(\edb_top_inst/n2584 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4118 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4119  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11] ), .O(\edb_top_inst/n2585 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4119 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4120  (.I0(\edb_top_inst/n2584 ), .I1(\edb_top_inst/n2583 ), 
            .I2(\edb_top_inst/n2585 ), .O(\edb_top_inst/n2586 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4120 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4121  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7] ), .O(\edb_top_inst/n2587 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4121 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4122  (.I0(\edb_top_inst/n2586 ), .I1(\edb_top_inst/n2587 ), 
            .O(\edb_top_inst/n2588 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4122 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4123  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6] ), 
            .I1(\edb_top_inst/n2582 ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I3(\edb_top_inst/n2588 ), .O(\edb_top_inst/n2589 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4123 .LUTMASK = 16'h7100;
    EFX_LUT4 \edb_top_inst/LUT__4124  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n2590 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4124 .LUTMASK = 16'h0b00;
    EFX_LUT4 \edb_top_inst/LUT__4125  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/n2591 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4125 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4126  (.I0(\edb_top_inst/n2590 ), .I1(\edb_top_inst/n2583 ), 
            .I2(\edb_top_inst/n2591 ), .I3(\edb_top_inst/n2586 ), .O(\edb_top_inst/n2592 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4126 .LUTMASK = 16'hbf00;
    EFX_LUT4 \edb_top_inst/LUT__4127  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/n2593 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4127 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4128  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/n2594 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4128 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4129  (.I0(\edb_top_inst/n2593 ), .I1(\edb_top_inst/n2594 ), 
            .O(\edb_top_inst/n2595 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4129 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4130  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13] ), .O(\edb_top_inst/n2596 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4130 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4131  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I2(\edb_top_inst/n2596 ), .O(\edb_top_inst/n2597 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4131 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__4132  (.I0(\edb_top_inst/n2592 ), .I1(\edb_top_inst/n2589 ), 
            .I2(\edb_top_inst/n2595 ), .I3(\edb_top_inst/n2597 ), .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4132 .LUTMASK = 16'hff10;
    EFX_LUT4 \edb_top_inst/LUT__4133  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n2598 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4133 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4134  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/n2599 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4134 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4135  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/n2600 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4135 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4136  (.I0(\edb_top_inst/n2598 ), .I1(\edb_top_inst/n2594 ), 
            .I2(\edb_top_inst/n2599 ), .I3(\edb_top_inst/n2600 ), .O(\edb_top_inst/n2601 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4136 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4137  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n2602 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4137 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4138  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/n2603 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4138 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4139  (.I0(\edb_top_inst/n2602 ), .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] ), .I3(\edb_top_inst/n2603 ), 
            .O(\edb_top_inst/n2604 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4139 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__4140  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n2605 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4140 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4141  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5] ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/n2606 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4141 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4142  (.I0(\edb_top_inst/n2601 ), .I1(\edb_top_inst/n2604 ), 
            .I2(\edb_top_inst/n2605 ), .I3(\edb_top_inst/n2606 ), .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/equal_9/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4142 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4143  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[8] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[15] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[15] ), 
            .O(\edb_top_inst/n2607 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4143 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4144  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[13] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[14] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[14] ), 
            .O(\edb_top_inst/n2608 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4144 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4145  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[11] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[12] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[12] ), 
            .O(\edb_top_inst/n2609 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4145 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4146  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[9] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[10] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[10] ), 
            .O(\edb_top_inst/n2610 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4146 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4147  (.I0(\edb_top_inst/n2607 ), .I1(\edb_top_inst/n2608 ), 
            .I2(\edb_top_inst/n2609 ), .I3(\edb_top_inst/n2610 ), .O(\edb_top_inst/n2611 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4147 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4148  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .O(\edb_top_inst/n2612 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4148 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4149  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .O(\edb_top_inst/n2613 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4149 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4150  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n2614 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4150 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4151  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .O(\edb_top_inst/n2615 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4151 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4152  (.I0(\edb_top_inst/n2612 ), .I1(\edb_top_inst/n2613 ), 
            .I2(\edb_top_inst/n2614 ), .I3(\edb_top_inst/n2615 ), .O(\edb_top_inst/n2616 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4152 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4153  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/n2611 ), .I3(\edb_top_inst/n2616 ), .O(\edb_top_inst/n2617 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haccc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4153 .LUTMASK = 16'haccc;
    EFX_LUT4 \edb_top_inst/LUT__4154  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n2618 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4154 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4155  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n2619 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4155 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__4156  (.I0(\edb_top_inst/n2618 ), .I1(\edb_top_inst/n2617 ), 
            .I2(\edb_top_inst/n2619 ), .I3(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n82 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f44, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4156 .LUTMASK = 16'h0f44;
    EFX_LUT4 \edb_top_inst/LUT__4157  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4157 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4158  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4158 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4159  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n69 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4159 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4160  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n68 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4160 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4161  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n67 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4161 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4162  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n66 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4162 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4163  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n65 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4163 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4164  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n64 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4164 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4165  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n63 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4165 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4166  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n62 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4166 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4167  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n61 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4167 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4168  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n60 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4168 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4169  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n59 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4169 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4170  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n58 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4170 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4171  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n57 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4171 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4172  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4172 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4173  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4173 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4174  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4174 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4175  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4175 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4176  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4176 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4177  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4177 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4178  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4178 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4179  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[8] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[8] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4179 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4180  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[9] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[9] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4180 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4181  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[10] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[10] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4181 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4182  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[11] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[11] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4182 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4183  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[12] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[12] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4183 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4184  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[13] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[13] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4184 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4185  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[14] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[14] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4185 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4186  (.I0(\edb_top_inst/la0/GEN_PROBE[3].this_probe_p1[15] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[15] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.trigger_cu/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4186 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4187  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4187 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4188  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4188 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4189  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), .O(\edb_top_inst/n2620 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4189 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4190  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n2621 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4190 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4191  (.I0(\edb_top_inst/n2620 ), .I1(\edb_top_inst/n2621 ), 
            .O(\edb_top_inst/n2622 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4191 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4192  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/n2623 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4192 .LUTMASK = 16'h8eaf;
    EFX_LUT4 \edb_top_inst/LUT__4193  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/n2622 ), .I3(\edb_top_inst/n2623 ), .O(\edb_top_inst/n2624 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4193 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4194  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/n2624 ), .O(\edb_top_inst/n2625 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4194 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__4195  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/n2625 ), .O(\edb_top_inst/n2626 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4195 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__4196  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7] ), 
            .I2(\edb_top_inst/n2626 ), .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4196 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__4197  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/n2627 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4197 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4198  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n2628 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4198 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4199  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n2629 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4199 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4200  (.I0(\edb_top_inst/n2621 ), .I1(\edb_top_inst/n2627 ), 
            .I2(\edb_top_inst/n2628 ), .I3(\edb_top_inst/n2629 ), .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4200 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4201  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n2630 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4201 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__4202  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n2631 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4202 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4203  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n2632 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4203 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4204  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n2633 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4204 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4205  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n2634 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4205 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4206  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n2635 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4206 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4207  (.I0(\edb_top_inst/n2632 ), .I1(\edb_top_inst/n2633 ), 
            .I2(\edb_top_inst/n2634 ), .I3(\edb_top_inst/n2635 ), .O(\edb_top_inst/n2636 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4207 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4208  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/n2631 ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n2636 ), .O(\edb_top_inst/n2637 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h752f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4208 .LUTMASK = 16'h752f;
    EFX_LUT4 \edb_top_inst/LUT__4209  (.I0(\edb_top_inst/n2637 ), .I1(\edb_top_inst/n2630 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[3].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4209 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4210  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4210 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4211  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4211 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4212  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4212 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4213  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4213 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4214  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4214 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4215  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4215 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4216  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[4].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4216 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4217  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4217 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4218  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4218 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4219  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4219 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4220  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4220 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4221  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4221 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4222  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4222 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4223  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[5].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.capture_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4223 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4224  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n40 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4224 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4225  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[0] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n22 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4225 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4226  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), .O(\edb_top_inst/n2638 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4226 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4227  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/n2639 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4227 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4228  (.I0(\edb_top_inst/n2638 ), .I1(\edb_top_inst/n2639 ), 
            .O(\edb_top_inst/n2640 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4228 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4229  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/n2641 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4229 .LUTMASK = 16'h8eaf;
    EFX_LUT4 \edb_top_inst/LUT__4230  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/n2640 ), .I3(\edb_top_inst/n2641 ), .O(\edb_top_inst/n2642 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4230 .LUTMASK = 16'hd4dd;
    EFX_LUT4 \edb_top_inst/LUT__4231  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/n2642 ), .O(\edb_top_inst/n2643 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4231 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__4232  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I2(\edb_top_inst/n2643 ), .O(\edb_top_inst/n2644 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4232 .LUTMASK = 16'hd4d4;
    EFX_LUT4 \edb_top_inst/LUT__4233  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I2(\edb_top_inst/n2644 ), .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n41 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4233 .LUTMASK = 16'h2b2b;
    EFX_LUT4 \edb_top_inst/LUT__4234  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/n2645 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4234 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4235  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/n2646 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4235 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4236  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] ), .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/n2647 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4236 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4237  (.I0(\edb_top_inst/n2639 ), .I1(\edb_top_inst/n2645 ), 
            .I2(\edb_top_inst/n2646 ), .I3(\edb_top_inst/n2647 ), .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/equal_9/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4237 .LUTMASK = 16'h7fff;
    EFX_LUT4 \edb_top_inst/LUT__4238  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .O(\edb_top_inst/n2648 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3dc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4238 .LUTMASK = 16'hc3dc;
    EFX_LUT4 \edb_top_inst/LUT__4239  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_gt ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp_eq ), 
            .O(\edb_top_inst/n2649 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4239 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4240  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[2] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[3] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[3] ), 
            .O(\edb_top_inst/n2650 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4240 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4241  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[4] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[5] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[5] ), 
            .O(\edb_top_inst/n2651 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4241 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4242  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[0] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[0] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[1] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[1] ), 
            .O(\edb_top_inst/n2652 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4242 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4243  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[6] ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp2[7] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/genblk1.genblk1.exp1[7] ), 
            .O(\edb_top_inst/n2653 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4243 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4244  (.I0(\edb_top_inst/n2650 ), .I1(\edb_top_inst/n2651 ), 
            .I2(\edb_top_inst/n2652 ), .I3(\edb_top_inst/n2653 ), .O(\edb_top_inst/n2654 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4244 .LUTMASK = 16'h8000;
    EFX_LUT4 \edb_top_inst/LUT__4245  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[0] ), 
            .I1(\edb_top_inst/n2649 ), .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[1] ), 
            .I3(\edb_top_inst/n2654 ), .O(\edb_top_inst/n2655 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h752f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4245 .LUTMASK = 16'h752f;
    EFX_LUT4 \edb_top_inst/LUT__4246  (.I0(\edb_top_inst/n2655 ), .I1(\edb_top_inst/n2648 ), 
            .I2(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[0].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n50 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4246 .LUTMASK = 16'h3535;
    EFX_LUT4 \edb_top_inst/LUT__4247  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n39 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4247 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4248  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n38 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4248 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4249  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n37 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4249 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4250  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n36 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4250 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4251  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n35 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4251 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4252  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4252 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4253  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[1].genblk1.internal_reg_pr[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4253 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4254  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[1] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[1] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n21 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4254 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4255  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[2] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n20 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4255 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4256  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[3] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n19 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4256 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4257  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[4] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[4] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n18 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4257 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4258  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[5] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[5] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n17 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4258 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4259  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[6] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[6] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n16 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4259 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4260  (.I0(\edb_top_inst/la0/GEN_PROBE[4].this_probe_p1[7] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[4].genblk7.GEN_REGS[2].genblk1.internal_reg_pr[7] ), 
            .O(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.trigger_cu/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4260 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4261  (.I0(\edb_top_inst/la0/la_trig_mask[1] ), 
            .I1(\edb_top_inst/la0/la_trig_mask[2] ), .I2(\edb_top_inst/la0/la_trig_mask[3] ), 
            .I3(\edb_top_inst/la0/la_trig_mask[4] ), .O(\edb_top_inst/n2656 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4261 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4262  (.I0(\edb_top_inst/la0/la_trig_mask[3] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[1] ), .I3(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n2657 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4262 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4263  (.I0(\edb_top_inst/la0/la_trig_mask[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I2(\edb_top_inst/la0/la_trig_mask[0] ), .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .O(\edb_top_inst/n2658 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4263 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4264  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[4] ), .I2(\edb_top_inst/n2657 ), 
            .I3(\edb_top_inst/n2658 ), .O(\edb_top_inst/n2659 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4264 .LUTMASK = 16'h7000;
    EFX_LUT4 \edb_top_inst/LUT__4265  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[2] ), .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[0] ), .O(\edb_top_inst/n2660 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4265 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4266  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[4] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk3.probe_cout ), 
            .I3(\edb_top_inst/la0/la_trig_mask[1] ), .O(\edb_top_inst/n2661 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4266 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4267  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk3.probe_cout ), 
            .I1(\edb_top_inst/la0/la_trig_mask[3] ), .I2(\edb_top_inst/n2660 ), 
            .I3(\edb_top_inst/n2661 ), .O(\edb_top_inst/n2662 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4267 .LUTMASK = 16'hb000;
    EFX_LUT4 \edb_top_inst/LUT__4268  (.I0(\edb_top_inst/n2659 ), .I1(\edb_top_inst/n2662 ), 
            .I2(\edb_top_inst/la0/la_trig_pattern[0] ), .I3(\edb_top_inst/la0/la_trig_pattern[1] ), 
            .O(\edb_top_inst/n2663 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha35c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4268 .LUTMASK = 16'ha35c;
    EFX_LUT4 \edb_top_inst/LUT__4269  (.I0(\edb_top_inst/n2656 ), .I1(\edb_top_inst/la0/la_trig_mask[0] ), 
            .I2(\edb_top_inst/n2663 ), .O(\edb_top_inst/la0/trigger_tu/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4269 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4270  (.I0(\edb_top_inst/la0/genblk2.la_capture_mask[1] ), 
            .I1(\edb_top_inst/la0/genblk2.la_capture_mask[2] ), .I2(\edb_top_inst/la0/genblk2.la_capture_mask[3] ), 
            .I3(\edb_top_inst/la0/genblk2.la_capture_mask[4] ), .O(\edb_top_inst/n2664 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4270 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4271  (.I0(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.cap_probe_cout ), 
            .I1(\edb_top_inst/la0/genblk2.la_capture_mask[3] ), .I2(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.cap_probe_cout ), 
            .I3(\edb_top_inst/la0/genblk2.la_capture_mask[1] ), .O(\edb_top_inst/n2665 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4271 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4272  (.I0(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.cap_probe_cout ), 
            .I1(\edb_top_inst/la0/genblk2.la_capture_mask[2] ), .I2(\edb_top_inst/la0/genblk2.la_capture_mask[0] ), 
            .I3(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.cap_probe_cout ), 
            .O(\edb_top_inst/n2666 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4272 .LUTMASK = 16'h0777;
    EFX_LUT4 \edb_top_inst/LUT__4273  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.cap_probe_cout ), 
            .I1(\edb_top_inst/la0/genblk2.la_capture_mask[4] ), .I2(\edb_top_inst/n2665 ), 
            .I3(\edb_top_inst/n2666 ), .O(\edb_top_inst/n2667 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4273 .LUTMASK = 16'h7000;
    EFX_LUT4 \edb_top_inst/LUT__4274  (.I0(\edb_top_inst/la0/GEN_PROBE[1].genblk7.genblk2.genblk1.cap_probe_cout ), 
            .I1(\edb_top_inst/la0/genblk2.la_capture_mask[1] ), .I2(\edb_top_inst/la0/GEN_PROBE[0].genblk7.genblk2.genblk1.cap_probe_cout ), 
            .I3(\edb_top_inst/la0/genblk2.la_capture_mask[0] ), .O(\edb_top_inst/n2668 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4274 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4275  (.I0(\edb_top_inst/la0/GEN_PROBE[4].genblk7.genblk2.genblk1.cap_probe_cout ), 
            .I1(\edb_top_inst/la0/genblk2.la_capture_mask[4] ), .I2(\edb_top_inst/la0/GEN_PROBE[3].genblk7.genblk2.genblk1.cap_probe_cout ), 
            .I3(\edb_top_inst/la0/genblk2.la_capture_mask[3] ), .O(\edb_top_inst/n2669 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4275 .LUTMASK = 16'hb0bb;
    EFX_LUT4 \edb_top_inst/LUT__4276  (.I0(\edb_top_inst/la0/genblk2.la_capture_mask[2] ), 
            .I1(\edb_top_inst/la0/GEN_PROBE[2].genblk7.genblk2.genblk1.cap_probe_cout ), 
            .I2(\edb_top_inst/n2668 ), .I3(\edb_top_inst/n2669 ), .O(\edb_top_inst/n2670 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4276 .LUTMASK = 16'hd000;
    EFX_LUT4 \edb_top_inst/LUT__4277  (.I0(\edb_top_inst/n2667 ), .I1(\edb_top_inst/n2670 ), 
            .I2(\edb_top_inst/la0/la_capture_pattern[0] ), .I3(\edb_top_inst/la0/la_capture_pattern[1] ), 
            .O(\edb_top_inst/n2671 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha35c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4277 .LUTMASK = 16'ha35c;
    EFX_LUT4 \edb_top_inst/LUT__4278  (.I0(\edb_top_inst/la0/genblk2.la_capture_mask[0] ), 
            .I1(\edb_top_inst/n2664 ), .I2(\edb_top_inst/n2671 ), .O(\edb_top_inst/la0/genblk2.global_capture_inst/n47 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4278 .LUTMASK = 16'hf4f4;
    EFX_LUT4 \edb_top_inst/LUT__4279  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n2672 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4279 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4280  (.I0(\edb_top_inst/n2672 ), .I1(\edb_top_inst/la0/la_window_depth[4] ), 
            .I2(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n2673 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4280 .LUTMASK = 16'hd3d3;
    EFX_LUT4 \edb_top_inst/LUT__4281  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I3(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n2674 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1ef1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4281 .LUTMASK = 16'h1ef1;
    EFX_LUT4 \edb_top_inst/LUT__4282  (.I0(\edb_top_inst/n2674 ), .I1(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I2(\edb_top_inst/la0/la_window_depth[3] ), .I3(\edb_top_inst/la0/la_trig_pos[8] ), 
            .O(\edb_top_inst/n2675 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h333a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4282 .LUTMASK = 16'h333a;
    EFX_LUT4 \edb_top_inst/LUT__4283  (.I0(\edb_top_inst/n2675 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/n2673 ), .I3(\edb_top_inst/la0/la_trig_pos[8] ), 
            .O(\edb_top_inst/n2676 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4114, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4283 .LUTMASK = 16'h4114;
    EFX_LUT4 \edb_top_inst/LUT__4284  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n2677 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4284 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4285  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n2678 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4285 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4286  (.I0(\edb_top_inst/n2677 ), .I1(\edb_top_inst/n2678 ), 
            .O(\edb_top_inst/n2679 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4286 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4287  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .I3(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n2680 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4287 .LUTMASK = 16'hf800;
    EFX_LUT4 \edb_top_inst/LUT__4288  (.I0(\edb_top_inst/n2672 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/n2680 ), 
            .O(\edb_top_inst/n2681 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4288 .LUTMASK = 16'h000d;
    EFX_LUT4 \edb_top_inst/LUT__4289  (.I0(\edb_top_inst/n2679 ), .I1(\edb_top_inst/n2681 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[11] ), .O(\edb_top_inst/n2682 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1e1e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4289 .LUTMASK = 16'h1e1e;
    EFX_LUT4 \edb_top_inst/LUT__4290  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n2683 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4290 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4291  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .I2(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I3(\edb_top_inst/n2683 ), .O(\edb_top_inst/n2684 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbffc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4291 .LUTMASK = 16'hbffc;
    EFX_LUT4 \edb_top_inst/LUT__4292  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[16] ), .O(\edb_top_inst/n2685 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heff0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4292 .LUTMASK = 16'heff0;
    EFX_LUT4 \edb_top_inst/LUT__4293  (.I0(\edb_top_inst/n2685 ), .I1(\edb_top_inst/la0/la_window_depth[4] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[9] ), .I3(\edb_top_inst/la0/la_window_depth[0] ), 
            .O(\edb_top_inst/n2686 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4293 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__4294  (.I0(\edb_top_inst/n2684 ), .I1(\edb_top_inst/la0/la_trig_pos[16] ), 
            .I2(\edb_top_inst/n2686 ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n2687 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4294 .LUTMASK = 16'h000e;
    EFX_LUT4 \edb_top_inst/LUT__4295  (.I0(\edb_top_inst/la0/la_trig_pos[16] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n2688 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4295 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__4296  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[9] ), .I2(\edb_top_inst/n2683 ), 
            .I3(\edb_top_inst/n2688 ), .O(\edb_top_inst/n2689 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4296 .LUTMASK = 16'h007d;
    EFX_LUT4 \edb_top_inst/LUT__4297  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n2690 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4297 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4298  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .I2(\edb_top_inst/la0/la_trig_pos[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .O(\edb_top_inst/n2691 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4298 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__4299  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/n2691 ), .O(\edb_top_inst/n2692 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4299 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4300  (.I0(\edb_top_inst/n2689 ), .I1(\edb_top_inst/n2690 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[7] ), .I3(\edb_top_inst/n2692 ), 
            .O(\edb_top_inst/n2693 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2c00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4300 .LUTMASK = 16'h2c00;
    EFX_LUT4 \edb_top_inst/LUT__4301  (.I0(\edb_top_inst/n2687 ), .I1(\edb_top_inst/n2682 ), 
            .I2(\edb_top_inst/n2676 ), .I3(\edb_top_inst/n2693 ), .O(\edb_top_inst/n2694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4301 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4302  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n2680 ), .O(\edb_top_inst/n2695 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4302 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4303  (.I0(\edb_top_inst/n2677 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[11] ), 
            .O(\edb_top_inst/n2696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4303 .LUTMASK = 16'h7878;
    EFX_LUT4 \edb_top_inst/LUT__4304  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I1(\edb_top_inst/n2696 ), .I2(\edb_top_inst/n2695 ), .O(\edb_top_inst/n2697 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4304 .LUTMASK = 16'he7e7;
    EFX_LUT4 \edb_top_inst/LUT__4305  (.I0(\edb_top_inst/n2672 ), .I1(\edb_top_inst/la0/la_window_depth[3] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n2698 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4305 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4306  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(\edb_top_inst/n2698 ), .O(\edb_top_inst/n2699 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4306 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4307  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/la0/la_window_depth[4] ), 
            .O(\edb_top_inst/n2700 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4307 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4308  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I3(\edb_top_inst/n2700 ), .O(\edb_top_inst/n2701 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hde3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4308 .LUTMASK = 16'hde3f;
    EFX_LUT4 \edb_top_inst/LUT__4309  (.I0(\edb_top_inst/n2677 ), .I1(\edb_top_inst/n2700 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), .O(\edb_top_inst/n2702 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4309 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__4310  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .I3(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n2703 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4310 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__4311  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(\edb_top_inst/n2703 ), .O(\edb_top_inst/n2704 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4311 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4312  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n2677 ), .I2(\edb_top_inst/n2690 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .O(\edb_top_inst/n2705 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4312 .LUTMASK = 16'h8f70;
    EFX_LUT4 \edb_top_inst/LUT__4313  (.I0(\edb_top_inst/n2701 ), .I1(\edb_top_inst/n2702 ), 
            .I2(\edb_top_inst/n2704 ), .I3(\edb_top_inst/n2705 ), .O(\edb_top_inst/n2706 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4313 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4314  (.I0(\edb_top_inst/n2672 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .I3(\edb_top_inst/n2690 ), 
            .O(\edb_top_inst/n2707 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4314 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__4315  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n2708 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4315 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4316  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n2708 ), .I2(\edb_top_inst/n2690 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .O(\edb_top_inst/n2709 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2fd0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4316 .LUTMASK = 16'h2fd0;
    EFX_LUT4 \edb_top_inst/LUT__4317  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/n2690 ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), .O(\edb_top_inst/n2710 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4317 .LUTMASK = 16'h8f70;
    EFX_LUT4 \edb_top_inst/LUT__4318  (.I0(\edb_top_inst/n2707 ), .I1(\edb_top_inst/n2709 ), 
            .I2(\edb_top_inst/n2710 ), .O(\edb_top_inst/n2711 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4318 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4319  (.I0(\edb_top_inst/n2697 ), .I1(\edb_top_inst/n2699 ), 
            .I2(\edb_top_inst/n2706 ), .I3(\edb_top_inst/n2711 ), .O(\edb_top_inst/n2712 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4319 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4320  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .O(\edb_top_inst/n2713 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4320 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4321  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/n2713 ), 
            .I3(\edb_top_inst/la0/la_trig_pos[13] ), .O(\edb_top_inst/n2714 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h40bf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4321 .LUTMASK = 16'h40bf;
    EFX_LUT4 \edb_top_inst/LUT__4322  (.I0(\edb_top_inst/n2708 ), .I1(\edb_top_inst/n2713 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .O(\edb_top_inst/n2715 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4322 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4323  (.I0(\edb_top_inst/n2677 ), .I1(\edb_top_inst/n2713 ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[14] ), 
            .O(\edb_top_inst/n2716 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h07f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4323 .LUTMASK = 16'h07f8;
    EFX_LUT4 \edb_top_inst/LUT__4324  (.I0(\edb_top_inst/n2716 ), .I1(\edb_top_inst/n2715 ), 
            .I2(\edb_top_inst/n2714 ), .I3(\edb_top_inst/la0/la_trig_pos[12] ), 
            .O(\edb_top_inst/n2717 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0140, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4324 .LUTMASK = 16'h0140;
    EFX_LUT4 \edb_top_inst/LUT__4325  (.I0(\edb_top_inst/n2680 ), .I1(\edb_top_inst/la0/la_trig_pos[15] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_trig_pos[10] ), 
            .O(\edb_top_inst/n2718 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dfe, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4325 .LUTMASK = 16'h3dfe;
    EFX_LUT4 \edb_top_inst/LUT__4326  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n2677 ), .I2(\edb_top_inst/n2690 ), .I3(\edb_top_inst/la0/la_trig_pos[6] ), 
            .O(\edb_top_inst/n2719 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h709f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4326 .LUTMASK = 16'h709f;
    EFX_LUT4 \edb_top_inst/LUT__4327  (.I0(\edb_top_inst/la0/la_trig_pos[6] ), 
            .I1(\edb_top_inst/n2700 ), .I2(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I3(\edb_top_inst/n2719 ), .O(\edb_top_inst/n2720 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4327 .LUTMASK = 16'hfb0f;
    EFX_LUT4 \edb_top_inst/LUT__4328  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/n2690 ), 
            .I3(\edb_top_inst/la0/la_trig_pos[5] ), .O(\edb_top_inst/n2721 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f70, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4328 .LUTMASK = 16'h8f70;
    EFX_LUT4 \edb_top_inst/LUT__4329  (.I0(\edb_top_inst/n2700 ), .I1(\edb_top_inst/la0/la_trig_pos[3] ), 
            .I2(\edb_top_inst/n2721 ), .O(\edb_top_inst/n2722 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4329 .LUTMASK = 16'h6060;
    EFX_LUT4 \edb_top_inst/LUT__4330  (.I0(\edb_top_inst/n2718 ), .I1(\edb_top_inst/n2720 ), 
            .I2(\edb_top_inst/n2717 ), .I3(\edb_top_inst/n2722 ), .O(\edb_top_inst/n2723 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4330 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4331  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I1(\edb_top_inst/n2696 ), .I2(\edb_top_inst/n2681 ), .O(\edb_top_inst/n2724 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7e7, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4331 .LUTMASK = 16'he7e7;
    EFX_LUT4 \edb_top_inst/LUT__4332  (.I0(\edb_top_inst/n2700 ), .I1(\edb_top_inst/la0/la_window_depth[0] ), 
            .I2(\edb_top_inst/la0/la_window_depth[1] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .O(\edb_top_inst/n2725 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd728, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4332 .LUTMASK = 16'hd728;
    EFX_LUT4 \edb_top_inst/LUT__4333  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/n2700 ), 
            .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), .O(\edb_top_inst/n2726 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4333 .LUTMASK = 16'hbf40;
    EFX_LUT4 \edb_top_inst/LUT__4334  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n2708 ), .I2(\edb_top_inst/n2690 ), .O(\edb_top_inst/n2727 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4334 .LUTMASK = 16'h9090;
    EFX_LUT4 \edb_top_inst/LUT__4335  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(\edb_top_inst/n2727 ), .I2(\edb_top_inst/n2725 ), .I3(\edb_top_inst/n2726 ), 
            .O(\edb_top_inst/n2728 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4335 .LUTMASK = 16'h6000;
    EFX_LUT4 \edb_top_inst/LUT__4336  (.I0(\edb_top_inst/n2708 ), .I1(\edb_top_inst/n2700 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), .O(\edb_top_inst/n2729 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4336 .LUTMASK = 16'hb4b4;
    EFX_LUT4 \edb_top_inst/LUT__4337  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_window_depth[3] ), .I2(\edb_top_inst/n2672 ), 
            .O(\edb_top_inst/n2730 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4337 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__4338  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(\edb_top_inst/n2730 ), .I2(\edb_top_inst/n2729 ), .O(\edb_top_inst/n2731 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4338 .LUTMASK = 16'h6060;
    EFX_LUT4 \edb_top_inst/LUT__4339  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I3(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n2732 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbcf1, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4339 .LUTMASK = 16'hbcf1;
    EFX_LUT4 \edb_top_inst/LUT__4340  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(\edb_top_inst/n2732 ), .I2(\edb_top_inst/n2690 ), .O(\edb_top_inst/n2733 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4340 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4341  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_window_depth[1] ), .I2(\edb_top_inst/la0/la_window_depth[2] ), 
            .O(\edb_top_inst/n2734 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e7e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4341 .LUTMASK = 16'h7e7e;
    EFX_LUT4 \edb_top_inst/LUT__4342  (.I0(\edb_top_inst/n2734 ), .I1(\edb_top_inst/n2690 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .O(\edb_top_inst/n2735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4342 .LUTMASK = 16'h7000;
    EFX_LUT4 \edb_top_inst/LUT__4343  (.I0(\edb_top_inst/la0/la_window_depth[3] ), 
            .I1(\edb_top_inst/n2672 ), .I2(\edb_top_inst/n2703 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .O(\edb_top_inst/n2736 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4fb0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4343 .LUTMASK = 16'h4fb0;
    EFX_LUT4 \edb_top_inst/LUT__4344  (.I0(\edb_top_inst/n2672 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), .I3(\edb_top_inst/n2690 ), 
            .O(\edb_top_inst/n2737 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ecf, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4344 .LUTMASK = 16'h7ecf;
    EFX_LUT4 \edb_top_inst/LUT__4345  (.I0(\edb_top_inst/n2735 ), .I1(\edb_top_inst/n2733 ), 
            .I2(\edb_top_inst/n2737 ), .I3(\edb_top_inst/n2736 ), .O(\edb_top_inst/n2738 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4345 .LUTMASK = 16'h0e00;
    EFX_LUT4 \edb_top_inst/LUT__4346  (.I0(\edb_top_inst/n2724 ), .I1(\edb_top_inst/n2728 ), 
            .I2(\edb_top_inst/n2731 ), .I3(\edb_top_inst/n2738 ), .O(\edb_top_inst/n2739 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4346 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4347  (.I0(\edb_top_inst/n2712 ), .I1(\edb_top_inst/n2723 ), 
            .I2(\edb_top_inst/n2694 ), .I3(\edb_top_inst/n2739 ), .O(\edb_top_inst/n2740 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4347 .LUTMASK = 16'h007f;
    EFX_LUT4 \edb_top_inst/LUT__4348  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .I2(\edb_top_inst/la0/la_trig_pos[2] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n2741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4348 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4349  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/la0/la_trig_pos[6] ), 
            .O(\edb_top_inst/n2742 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4349 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4350  (.I0(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[8] ), .I2(\edb_top_inst/n2741 ), 
            .I3(\edb_top_inst/n2742 ), .O(\edb_top_inst/n2743 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4350 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4351  (.I0(\edb_top_inst/la0/la_trig_pos[12] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[13] ), .I2(\edb_top_inst/la0/la_trig_pos[14] ), 
            .I3(\edb_top_inst/la0/la_trig_pos[15] ), .O(\edb_top_inst/n2744 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4351 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4352  (.I0(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[16] ), .I2(\edb_top_inst/n2744 ), 
            .O(\edb_top_inst/n2745 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4352 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4353  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[10] ), .I2(\edb_top_inst/n2743 ), 
            .I3(\edb_top_inst/n2745 ), .O(\edb_top_inst/n2746 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4353 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4354  (.I0(\edb_top_inst/la0/la_num_trigger[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), .O(\edb_top_inst/n2747 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4354 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4355  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .I2(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[3] ), .O(\edb_top_inst/n2748 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4355 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4356  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[5] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I3(\edb_top_inst/n2748 ), .O(\edb_top_inst/n2749 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4356 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4357  (.I0(\edb_top_inst/la0/la_num_trigger[6] ), 
            .I1(\edb_top_inst/n2747 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I3(\edb_top_inst/n2749 ), .O(\edb_top_inst/n2750 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4200, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4357 .LUTMASK = 16'h4200;
    EFX_LUT4 \edb_top_inst/LUT__4358  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/n2748 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[5] ), .O(\edb_top_inst/n2751 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4bf4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4358 .LUTMASK = 16'h4bf4;
    EFX_LUT4 \edb_top_inst/LUT__4359  (.I0(\edb_top_inst/n2747 ), .I1(\edb_top_inst/n2751 ), 
            .I2(\edb_top_inst/la0/la_num_trigger[6] ), .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .O(\edb_top_inst/n2752 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4359 .LUTMASK = 16'h1001;
    EFX_LUT4 \edb_top_inst/LUT__4360  (.I0(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[9] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .O(\edb_top_inst/n2753 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4360 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__4361  (.I0(\edb_top_inst/la0/la_num_trigger[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .I2(\edb_top_inst/la0/la_num_trigger[9] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), .O(\edb_top_inst/n2754 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4361 .LUTMASK = 16'h9009;
    EFX_LUT4 \edb_top_inst/LUT__4362  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[5] ), .I2(\edb_top_inst/la0/la_num_trigger[6] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[7] ), .O(\edb_top_inst/n2755 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4362 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4363  (.I0(\edb_top_inst/n2753 ), .I1(\edb_top_inst/n2754 ), 
            .I2(\edb_top_inst/n2748 ), .I3(\edb_top_inst/n2755 ), .O(\edb_top_inst/n2756 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ccc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4363 .LUTMASK = 16'h5ccc;
    EFX_LUT4 \edb_top_inst/LUT__4364  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .O(\edb_top_inst/n2757 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4364 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4365  (.I0(\edb_top_inst/la0/la_num_trigger[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .O(\edb_top_inst/n2758 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4365 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4366  (.I0(\edb_top_inst/la0/la_num_trigger[2] ), 
            .I1(\edb_top_inst/n2758 ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I3(\edb_top_inst/n2757 ), .O(\edb_top_inst/n2759 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdde, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4366 .LUTMASK = 16'hbdde;
    EFX_LUT4 \edb_top_inst/LUT__4367  (.I0(\edb_top_inst/la0/la_num_trigger[0] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[1] ), .I2(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .O(\edb_top_inst/n2760 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb7d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4367 .LUTMASK = 16'heb7d;
    EFX_LUT4 \edb_top_inst/LUT__4368  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), .O(\edb_top_inst/n2761 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4368 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4369  (.I0(\edb_top_inst/la0/la_num_trigger[14] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[15] ), .I2(\edb_top_inst/la0/la_num_trigger[16] ), 
            .O(\edb_top_inst/n2762 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4369 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4370  (.I0(\edb_top_inst/la0/la_num_trigger[12] ), 
            .I1(\edb_top_inst/n2748 ), .I2(\edb_top_inst/n2761 ), .I3(\edb_top_inst/n2762 ), 
            .O(\edb_top_inst/n2763 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4370 .LUTMASK = 16'h4100;
    EFX_LUT4 \edb_top_inst/LUT__4371  (.I0(\edb_top_inst/n2759 ), .I1(\edb_top_inst/n2760 ), 
            .I2(\edb_top_inst/n2756 ), .I3(\edb_top_inst/n2763 ), .O(\edb_top_inst/n2764 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4371 .LUTMASK = 16'h1000;
    EFX_LUT4 \edb_top_inst/LUT__4372  (.I0(\edb_top_inst/la0/la_num_trigger[5] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[6] ), .I2(\edb_top_inst/la0/la_num_trigger[7] ), 
            .O(\edb_top_inst/n2765 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4372 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4373  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[8] ), .I2(\edb_top_inst/la0/la_num_trigger[9] ), 
            .I3(\edb_top_inst/la0/la_num_trigger[10] ), .O(\edb_top_inst/n2766 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4373 .LUTMASK = 16'h0001;
    EFX_LUT4 \edb_top_inst/LUT__4374  (.I0(\edb_top_inst/n2748 ), .I1(\edb_top_inst/n2765 ), 
            .I2(\edb_top_inst/n2766 ), .O(\edb_top_inst/n2767 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4374 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4375  (.I0(\edb_top_inst/la0/la_num_trigger[4] ), 
            .I1(\edb_top_inst/la0/la_num_trigger[8] ), .I2(\edb_top_inst/la0/la_num_trigger[9] ), 
            .O(\edb_top_inst/n2768 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4375 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4376  (.I0(\edb_top_inst/la0/la_num_trigger[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), .O(\edb_top_inst/n2769 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4376 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4377  (.I0(\edb_top_inst/n2748 ), .I1(\edb_top_inst/n2765 ), 
            .I2(\edb_top_inst/n2768 ), .I3(\edb_top_inst/n2769 ), .O(\edb_top_inst/n2770 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4377 .LUTMASK = 16'h7f80;
    EFX_LUT4 \edb_top_inst/LUT__4378  (.I0(\edb_top_inst/la0/la_num_trigger[13] ), 
            .I1(\edb_top_inst/n2770 ), .I2(\edb_top_inst/n2767 ), .I3(\edb_top_inst/la0/la_num_trigger[11] ), 
            .O(\edb_top_inst/n2771 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4378 .LUTMASK = 16'h1001;
    EFX_LUT4 \edb_top_inst/LUT__4379  (.I0(\edb_top_inst/n2752 ), .I1(\edb_top_inst/n2750 ), 
            .I2(\edb_top_inst/n2764 ), .I3(\edb_top_inst/n2771 ), .O(\edb_top_inst/n2772 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4379 .LUTMASK = 16'he000;
    EFX_LUT4 \edb_top_inst/LUT__4380  (.I0(\edb_top_inst/n2746 ), .I1(\edb_top_inst/n2772 ), 
            .O(\edb_top_inst/n2773 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4380 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4381  (.I0(\edb_top_inst/n2740 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I2(\edb_top_inst/n2773 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n2774 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4381 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4382  (.I0(\edb_top_inst/la0/tu_trigger ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n2775 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4382 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4383  (.I0(\edb_top_inst/la0/la_biu_inst/run_trig_p2 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/run_trig_imdt_p2 ), .O(\edb_top_inst/n2776 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4383 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4384  (.I0(\edb_top_inst/n2746 ), .I1(\edb_top_inst/n2776 ), 
            .I2(\edb_top_inst/n2775 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n2777 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4384 .LUTMASK = 16'hf0ee;
    EFX_LUT4 \edb_top_inst/LUT__4385  (.I0(\edb_top_inst/la0/la_trig_pos[8] ), 
            .I1(\edb_top_inst/n2698 ), .O(\edb_top_inst/n2778 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4385 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4386  (.I0(\edb_top_inst/n2672 ), .I1(\edb_top_inst/la0/la_trig_pos[7] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[0] ), .I3(\edb_top_inst/n2690 ), 
            .O(\edb_top_inst/n2779 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hed3f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4386 .LUTMASK = 16'hed3f;
    EFX_LUT4 \edb_top_inst/LUT__4387  (.I0(\edb_top_inst/la0/la_window_depth[2] ), 
            .I1(\edb_top_inst/n2708 ), .I2(\edb_top_inst/n2690 ), .I3(\edb_top_inst/la0/la_trig_pos[4] ), 
            .O(\edb_top_inst/n2780 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2fd0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4387 .LUTMASK = 16'h2fd0;
    EFX_LUT4 \edb_top_inst/LUT__4388  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n2781 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4388 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4389  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_window_depth[0] ), .I2(\edb_top_inst/n2781 ), 
            .I3(\edb_top_inst/la0/la_trig_pos[16] ), .O(\edb_top_inst/n2782 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f8a, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4389 .LUTMASK = 16'h7f8a;
    EFX_LUT4 \edb_top_inst/LUT__4390  (.I0(\edb_top_inst/n2695 ), .I1(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I2(\edb_top_inst/n2782 ), .I3(\edb_top_inst/n2780 ), .O(\edb_top_inst/n2783 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4390 .LUTMASK = 16'h0700;
    EFX_LUT4 \edb_top_inst/LUT__4391  (.I0(\edb_top_inst/n2683 ), .I1(\edb_top_inst/n2690 ), 
            .I2(\edb_top_inst/la0/la_trig_pos[1] ), .O(\edb_top_inst/n2784 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4391 .LUTMASK = 16'h7878;
    EFX_LUT4 \edb_top_inst/LUT__4392  (.I0(\edb_top_inst/n2690 ), .I1(\edb_top_inst/la0/la_trig_pos[11] ), 
            .I2(\edb_top_inst/n2678 ), .O(\edb_top_inst/n2785 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4392 .LUTMASK = 16'h3e3e;
    EFX_LUT4 \edb_top_inst/LUT__4393  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/n2703 ), .I2(\edb_top_inst/n2784 ), .I3(\edb_top_inst/n2785 ), 
            .O(\edb_top_inst/n2786 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4393 .LUTMASK = 16'h6000;
    EFX_LUT4 \edb_top_inst/LUT__4394  (.I0(\edb_top_inst/n2779 ), .I1(\edb_top_inst/n2778 ), 
            .I2(\edb_top_inst/n2783 ), .I3(\edb_top_inst/n2786 ), .O(\edb_top_inst/n2787 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4394 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4395  (.I0(\edb_top_inst/n2787 ), .I1(\edb_top_inst/n2723 ), 
            .I2(\edb_top_inst/n2777 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n2788 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf70f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4395 .LUTMASK = 16'hf70f;
    EFX_LUT4 \edb_top_inst/LUT__4396  (.I0(\edb_top_inst/la0/la_stop_trig ), 
            .I1(\edb_top_inst/n2775 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n2789 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4396 .LUTMASK = 16'hf400;
    EFX_LUT4 \edb_top_inst/LUT__4397  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[10] ), .O(\edb_top_inst/n2790 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4397 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4398  (.I0(\edb_top_inst/n2790 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[9] ), .I3(\edb_top_inst/n2743 ), 
            .O(\edb_top_inst/n2791 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4398 .LUTMASK = 16'he7be;
    EFX_LUT4 \edb_top_inst/LUT__4399  (.I0(\edb_top_inst/n2741 ), .I1(\edb_top_inst/n2742 ), 
            .O(\edb_top_inst/n2792 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4399 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4400  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[8] ), .O(\edb_top_inst/n2793 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4400 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4401  (.I0(\edb_top_inst/n2793 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[7] ), .I3(\edb_top_inst/n2792 ), 
            .O(\edb_top_inst/n2794 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4401 .LUTMASK = 16'he7be;
    EFX_LUT4 \edb_top_inst/LUT__4402  (.I0(\edb_top_inst/la0/la_trig_pos[9] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[10] ), .I2(\edb_top_inst/n2743 ), 
            .I3(\edb_top_inst/la0/la_trig_pos[11] ), .O(\edb_top_inst/n2795 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4402 .LUTMASK = 16'hef10;
    EFX_LUT4 \edb_top_inst/LUT__4403  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .O(\edb_top_inst/n2796 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4403 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4404  (.I0(\edb_top_inst/n2796 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[4] ), .I3(\edb_top_inst/n2741 ), 
            .O(\edb_top_inst/n2797 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4404 .LUTMASK = 16'he7be;
    EFX_LUT4 \edb_top_inst/LUT__4405  (.I0(\edb_top_inst/la0/la_trig_pos[0] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[1] ), .O(\edb_top_inst/n2798 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4405 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4406  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[3] ), .O(\edb_top_inst/n2799 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4406 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4407  (.I0(\edb_top_inst/n2799 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I2(\edb_top_inst/la0/la_trig_pos[2] ), .I3(\edb_top_inst/n2798 ), 
            .O(\edb_top_inst/n2800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he7be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4407 .LUTMASK = 16'he7be;
    EFX_LUT4 \edb_top_inst/LUT__4408  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[6] ), .O(\edb_top_inst/n2801 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4408 .LUTMASK = 16'h6666;
    EFX_LUT4 \edb_top_inst/LUT__4409  (.I0(\edb_top_inst/la0/la_trig_pos[4] ), 
            .I1(\edb_top_inst/la0/la_trig_pos[5] ), .I2(\edb_top_inst/n2741 ), 
            .I3(\edb_top_inst/n2801 ), .O(\edb_top_inst/n2802 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef10, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4409 .LUTMASK = 16'hef10;
    EFX_LUT4 \edb_top_inst/LUT__4410  (.I0(\edb_top_inst/la0/la_trig_pos[16] ), 
            .I1(\edb_top_inst/n2691 ), .I2(\edb_top_inst/n2744 ), .O(\edb_top_inst/n2803 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4410 .LUTMASK = 16'h1010;
    EFX_LUT4 \edb_top_inst/LUT__4411  (.I0(\edb_top_inst/n2797 ), .I1(\edb_top_inst/n2800 ), 
            .I2(\edb_top_inst/n2802 ), .I3(\edb_top_inst/n2803 ), .O(\edb_top_inst/n2804 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4411 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4412  (.I0(\edb_top_inst/n2791 ), .I1(\edb_top_inst/n2794 ), 
            .I2(\edb_top_inst/n2795 ), .I3(\edb_top_inst/n2804 ), .O(\edb_top_inst/n2805 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4412 .LUTMASK = 16'h0100;
    EFX_LUT4 \edb_top_inst/LUT__4413  (.I0(\edb_top_inst/n2805 ), .I1(\edb_top_inst/n2789 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n2806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d03, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4413 .LUTMASK = 16'h0d03;
    EFX_LUT4 \edb_top_inst/LUT__4414  (.I0(\edb_top_inst/n2788 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I2(\edb_top_inst/n2806 ), .O(\edb_top_inst/n2807 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4414 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__4415  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n2805 ), .O(\edb_top_inst/n2808 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4415 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4416  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n2809 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4416 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4417  (.I0(\edb_top_inst/n2808 ), .I1(\edb_top_inst/n2809 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/n2810 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4417 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4418  (.I0(\edb_top_inst/n2775 ), .I1(\edb_top_inst/n2712 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n2811 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4418 .LUTMASK = 16'h0a0c;
    EFX_LUT4 \edb_top_inst/LUT__4419  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/n2811 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .O(\edb_top_inst/n2812 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4419 .LUTMASK = 16'hd0d0;
    EFX_LUT4 \edb_top_inst/LUT__4420  (.I0(\edb_top_inst/n2774 ), .I1(\edb_top_inst/n2807 ), 
            .I2(\edb_top_inst/n2810 ), .I3(\edb_top_inst/n2812 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4420 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__4421  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .O(\edb_top_inst/n2813 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05fc, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4421 .LUTMASK = 16'h05fc;
    EFX_LUT4 \edb_top_inst/LUT__4422  (.I0(\edb_top_inst/la0/la_stop_trig ), 
            .I1(\edb_top_inst/la0/capture_enable ), .I2(\edb_top_inst/n2813 ), 
            .O(\edb_top_inst/la0/la_biu_inst/n1182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4422 .LUTMASK = 16'hefef;
    EFX_LUT4 \edb_top_inst/LUT__4423  (.I0(\edb_top_inst/n2360 ), .I1(\edb_top_inst/la0/biu_ready ), 
            .O(\edb_top_inst/la0/la_biu_inst/n369 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4423 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4424  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), .O(\edb_top_inst/la0/la_biu_inst/n1285 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4424 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4425  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2 ), .I2(\edb_top_inst/la0/la_biu_inst/str_sync_wbff2q ), 
            .I3(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00be, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4425 .LUTMASK = 16'h00be;
    EFX_LUT4 \edb_top_inst/LUT__4426  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), 
            .I1(\edb_top_inst/la0/la_resetn ), .I2(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .O(\edb_top_inst/ceg_net351 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4426 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4427  (.I0(\edb_top_inst/n2775 ), .I1(\edb_top_inst/n2787 ), 
            .I2(\edb_top_inst/n2723 ), .O(\edb_top_inst/n2814 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4427 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4428  (.I0(\edb_top_inst/n2740 ), .I1(\edb_top_inst/n2773 ), 
            .I2(\edb_top_inst/n2814 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n2815 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4428 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4429  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .O(\edb_top_inst/n2816 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4429 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4430  (.I0(\edb_top_inst/n2775 ), .I1(\edb_top_inst/n2772 ), 
            .I2(\edb_top_inst/n2712 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n2817 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hee0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4430 .LUTMASK = 16'hee0f;
    EFX_LUT4 \edb_top_inst/LUT__4431  (.I0(\edb_top_inst/n2817 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .O(\edb_top_inst/n2818 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4431 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4432  (.I0(\edb_top_inst/n2815 ), .I1(\edb_top_inst/n2816 ), 
            .I2(\edb_top_inst/n2818 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .O(\edb_top_inst/la0/la_biu_inst/next_state[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4432 .LUTMASK = 16'h00f4;
    EFX_LUT4 \edb_top_inst/LUT__4433  (.I0(\edb_top_inst/n2772 ), .I1(\edb_top_inst/n2746 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .O(\edb_top_inst/n2819 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4433 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__4434  (.I0(\edb_top_inst/n2787 ), .I1(\edb_top_inst/n2723 ), 
            .I2(\edb_top_inst/n2772 ), .I3(\edb_top_inst/n2775 ), .O(\edb_top_inst/n2820 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4434 .LUTMASK = 16'h008f;
    EFX_LUT4 \edb_top_inst/LUT__4435  (.I0(\edb_top_inst/n2775 ), .I1(\edb_top_inst/la0/la_stop_trig ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .O(\edb_top_inst/n2821 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4435 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4436  (.I0(\edb_top_inst/n2740 ), .I1(\edb_top_inst/n2819 ), 
            .I2(\edb_top_inst/n2820 ), .I3(\edb_top_inst/n2821 ), .O(\edb_top_inst/n2822 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4436 .LUTMASK = 16'hf0bb;
    EFX_LUT4 \edb_top_inst/LUT__4437  (.I0(\edb_top_inst/n2775 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .O(\edb_top_inst/n2823 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4437 .LUTMASK = 16'h4040;
    EFX_LUT4 \edb_top_inst/LUT__4438  (.I0(\edb_top_inst/n2772 ), .I1(\edb_top_inst/n2823 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), .I3(\edb_top_inst/n2712 ), 
            .O(\edb_top_inst/n2824 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7770, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4438 .LUTMASK = 16'h7770;
    EFX_LUT4 \edb_top_inst/LUT__4439  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n2825 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0140, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4439 .LUTMASK = 16'h0140;
    EFX_LUT4 \edb_top_inst/LUT__4440  (.I0(\edb_top_inst/n2824 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .I3(\edb_top_inst/n2825 ), 
            .O(\edb_top_inst/n2826 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4440 .LUTMASK = 16'h00ef;
    EFX_LUT4 \edb_top_inst/LUT__4441  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n2822 ), .I2(\edb_top_inst/n2816 ), .I3(\edb_top_inst/n2826 ), 
            .O(\edb_top_inst/la0/la_biu_inst/next_state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h10ff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4441 .LUTMASK = 16'h10ff;
    EFX_LUT4 \edb_top_inst/LUT__4442  (.I0(\edb_top_inst/n2723 ), .I1(\edb_top_inst/n2787 ), 
            .I2(\edb_top_inst/n2772 ), .O(\edb_top_inst/n2827 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4442 .LUTMASK = 16'h7878;
    EFX_LUT4 \edb_top_inst/LUT__4443  (.I0(\edb_top_inst/n2827 ), .I1(\edb_top_inst/n2775 ), 
            .I2(\edb_top_inst/n2821 ), .O(\edb_top_inst/n2828 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4443 .LUTMASK = 16'he0e0;
    EFX_LUT4 \edb_top_inst/LUT__4444  (.I0(\edb_top_inst/n2772 ), .I1(\edb_top_inst/n2746 ), 
            .O(\edb_top_inst/n2829 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4444 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4445  (.I0(\edb_top_inst/n2740 ), .I1(\edb_top_inst/n2829 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .O(\edb_top_inst/n2830 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4445 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__4446  (.I0(\edb_top_inst/n2776 ), .I1(\edb_top_inst/n2746 ), 
            .O(\edb_top_inst/n2831 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4446 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4447  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I1(\edb_top_inst/n2805 ), .I2(\edb_top_inst/n2831 ), .I3(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .O(\edb_top_inst/n2832 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4447 .LUTMASK = 16'heef8;
    EFX_LUT4 \edb_top_inst/LUT__4448  (.I0(\edb_top_inst/n2832 ), .I1(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n2833 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4448 .LUTMASK = 16'h0d0d;
    EFX_LUT4 \edb_top_inst/LUT__4449  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[1] ), 
            .I1(\edb_top_inst/n2805 ), .I2(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), 
            .I3(\edb_top_inst/la0/la_biu_inst/curr_state[2] ), .O(\edb_top_inst/n2834 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4449 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__4450  (.I0(\edb_top_inst/n2809 ), .I1(\edb_top_inst/n2811 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), .I3(\edb_top_inst/n2834 ), 
            .O(\edb_top_inst/n2835 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4450 .LUTMASK = 16'h001f;
    EFX_LUT4 \edb_top_inst/LUT__4451  (.I0(\edb_top_inst/n2828 ), .I1(\edb_top_inst/n2830 ), 
            .I2(\edb_top_inst/n2833 ), .I3(\edb_top_inst/n2835 ), .O(\edb_top_inst/la0/la_biu_inst/next_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4451 .LUTMASK = 16'h004f;
    EFX_LUT4 \edb_top_inst/LUT__4452  (.I0(\edb_top_inst/la0/la_biu_inst/n369 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2q ), .I2(\edb_top_inst/la0/la_biu_inst/rdy_sync_tff2 ), 
            .O(\edb_top_inst/ceg_net348 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4452 .LUTMASK = 16'h4141;
    EFX_LUT4 \edb_top_inst/LUT__4453  (.I0(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/axi_fsm_state[0] ), .O(\edb_top_inst/la0/la_biu_inst/next_fsm_state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4453 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4454  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/n2816 ), 
            .I3(\edb_top_inst/n2775 ), .O(\edb_top_inst/la0/la_biu_inst/n2027 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefff, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4454 .LUTMASK = 16'hefff;
    EFX_LUT4 \edb_top_inst/LUT__4455  (.I0(\edb_top_inst/n2813 ), .I1(\edb_top_inst/la0/capture_enable ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_push )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4455 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4456  (.I0(\edb_top_inst/la0/la_biu_inst/n2027 ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_push ), .O(\edb_top_inst/n2836 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4456 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4457  (.I0(\edb_top_inst/n2712 ), .I1(\edb_top_inst/n2836 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4457 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4458  (.I0(\edb_top_inst/la0/la_biu_inst/curr_state[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/curr_state[3] ), .I2(\edb_top_inst/n2809 ), 
            .I3(\edb_top_inst/la0/la_resetn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_rstn )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4458 .LUTMASK = 16'hef00;
    EFX_LUT4 \edb_top_inst/LUT__4459  (.I0(\edb_top_inst/la0/la_biu_inst/n2027 ), 
            .I1(\edb_top_inst/la0/capture_enable ), .O(\edb_top_inst/la0/la_biu_inst/fifo_pop )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4459 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4460  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/is_last_data ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n800 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4460 .LUTMASK = 16'hbbbb;
    EFX_LUT4 \edb_top_inst/LUT__4461  (.I0(\edb_top_inst/n2836 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_rstn ), 
            .O(\edb_top_inst/ceg_net355 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4461 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4462  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/pop_p2 ), 
            .I1(\edb_top_inst/n2417 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4462 .LUTMASK = 16'heeee;
    EFX_LUT4 \edb_top_inst/LUT__4463  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[15] ), .I2(\edb_top_inst/n2417 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4463 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4464  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[16] ), .I2(\edb_top_inst/n2417 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4464 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4465  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[17] ), .I2(\edb_top_inst/n2417 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4465 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4466  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[18] ), .I2(\edb_top_inst/n2417 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4466 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4467  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[19] ), .I2(\edb_top_inst/n2417 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4467 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4468  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[20] ), .I2(\edb_top_inst/n2417 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4468 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4469  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[21] ), .I2(\edb_top_inst/n2417 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4469 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4470  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[22] ), .I2(\edb_top_inst/n2417 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4470 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4471  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[23] ), .I2(\edb_top_inst/n2417 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4471 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4472  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[24] ), .I2(\edb_top_inst/n2417 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4472 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4473  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/rd_pointer[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/addr_reg[25] ), .I2(\edb_top_inst/n2417 ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4473 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4474  (.I0(\edb_top_inst/n2679 ), .I1(\edb_top_inst/n2681 ), 
            .O(\edb_top_inst/n2837 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4474 .LUTMASK = 16'h1111;
    EFX_LUT4 \edb_top_inst/LUT__4475  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I1(\edb_top_inst/n2708 ), .O(\edb_top_inst/n2838 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4475 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4476  (.I0(\edb_top_inst/n2700 ), .I1(\edb_top_inst/n2838 ), 
            .I2(\edb_top_inst/n2837 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4476 .LUTMASK = 16'h8f88;
    EFX_LUT4 \edb_top_inst/LUT__4477  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/n2713 ), .I2(\edb_top_inst/n2781 ), .O(\edb_top_inst/n2839 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4477 .LUTMASK = 16'h0101;
    EFX_LUT4 \edb_top_inst/LUT__4478  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .O(\edb_top_inst/n2840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4478 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4479  (.I0(\edb_top_inst/n2840 ), .I1(\edb_top_inst/n2690 ), 
            .I2(\edb_top_inst/n2683 ), .O(\edb_top_inst/n2841 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4479 .LUTMASK = 16'h8080;
    EFX_LUT4 \edb_top_inst/LUT__4480  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I1(\edb_top_inst/n2839 ), .I2(\edb_top_inst/n2841 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4480 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4481  (.I0(\edb_top_inst/n2677 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n2842 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030e, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4481 .LUTMASK = 16'h030e;
    EFX_LUT4 \edb_top_inst/LUT__4482  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .O(\edb_top_inst/n2843 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4482 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4483  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .I2(\edb_top_inst/n2843 ), 
            .I3(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n2844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4483 .LUTMASK = 16'hbb0f;
    EFX_LUT4 \edb_top_inst/LUT__4484  (.I0(\edb_top_inst/n2844 ), .I1(\edb_top_inst/n2700 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .I3(\edb_top_inst/n2842 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4484 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4485  (.I0(\edb_top_inst/la0/la_window_depth[4] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .I2(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n2845 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4485 .LUTMASK = 16'h1414;
    EFX_LUT4 \edb_top_inst/LUT__4486  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .O(\edb_top_inst/n2846 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4486 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4487  (.I0(\edb_top_inst/n2846 ), .I1(\edb_top_inst/n2840 ), 
            .I2(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n2847 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4487 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4488  (.I0(\edb_top_inst/n2847 ), .I1(\edb_top_inst/n2700 ), 
            .O(\edb_top_inst/n2848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4488 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4489  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I1(\edb_top_inst/n2845 ), .I2(\edb_top_inst/n2848 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4489 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4490  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n2849 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4490 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4491  (.I0(\edb_top_inst/la0/la_window_depth[0] ), 
            .I1(\edb_top_inst/n2849 ), .O(\edb_top_inst/n2850 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4491 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4492  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .I2(\edb_top_inst/la0/la_window_depth[0] ), 
            .O(\edb_top_inst/n2851 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4492 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4493  (.I0(\edb_top_inst/n2851 ), .I1(\edb_top_inst/n2843 ), 
            .I2(\edb_top_inst/la0/la_window_depth[1] ), .O(\edb_top_inst/n2852 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4493 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4494  (.I0(\edb_top_inst/n2852 ), .I1(\edb_top_inst/n2838 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n2690 ), 
            .O(\edb_top_inst/n2853 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4494 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4495  (.I0(\edb_top_inst/n2850 ), .I1(\edb_top_inst/n2845 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I3(\edb_top_inst/n2853 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4495 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4496  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/n2840 ), .O(\edb_top_inst/n2854 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4496 .LUTMASK = 16'h4444;
    EFX_LUT4 \edb_top_inst/LUT__4497  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2855 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4497 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4498  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2856 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4498 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4499  (.I0(\edb_top_inst/n2856 ), .I1(\edb_top_inst/n2855 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2857 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4499 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4500  (.I0(\edb_top_inst/n2857 ), .I1(\edb_top_inst/n2854 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n2690 ), 
            .O(\edb_top_inst/n2858 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4500 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4501  (.I0(\edb_top_inst/n2849 ), .I1(\edb_top_inst/n2845 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I3(\edb_top_inst/n2858 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4501 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4502  (.I0(\edb_top_inst/n2677 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/n2845 ), .O(\edb_top_inst/n2859 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4502 .LUTMASK = 16'hb0b0;
    EFX_LUT4 \edb_top_inst/LUT__4503  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2860 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4503 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4504  (.I0(\edb_top_inst/n2860 ), .I1(\edb_top_inst/n2856 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2861 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4504 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4505  (.I0(\edb_top_inst/n2861 ), .I1(\edb_top_inst/n2844 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n2690 ), 
            .O(\edb_top_inst/n2862 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4505 .LUTMASK = 16'h3a00;
    EFX_LUT4 \edb_top_inst/LUT__4506  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I1(\edb_top_inst/n2859 ), .I2(\edb_top_inst/n2862 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4506 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4507  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2863 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4507 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4508  (.I0(\edb_top_inst/n2863 ), .I1(\edb_top_inst/n2860 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2864 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4508 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4509  (.I0(\edb_top_inst/n2864 ), .I1(\edb_top_inst/n2847 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n2690 ), 
            .O(\edb_top_inst/n2865 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4509 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4510  (.I0(\edb_top_inst/n2678 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I2(\edb_top_inst/n2865 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4510 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4511  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2866 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4511 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4512  (.I0(\edb_top_inst/n2866 ), .I1(\edb_top_inst/n2863 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2867 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4512 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4513  (.I0(\edb_top_inst/n2867 ), .I1(\edb_top_inst/n2852 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .O(\edb_top_inst/n2868 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4513 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4514  (.I0(\edb_top_inst/n2868 ), .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), 
            .I2(\edb_top_inst/la0/la_window_depth[3] ), .I3(\edb_top_inst/n2698 ), 
            .O(\edb_top_inst/n2869 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4514 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4515  (.I0(\edb_top_inst/n2708 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I3(\edb_top_inst/n2869 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4515 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4516  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2870 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4516 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4517  (.I0(\edb_top_inst/n2870 ), .I1(\edb_top_inst/n2866 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2871 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4517 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4518  (.I0(\edb_top_inst/n2871 ), .I1(\edb_top_inst/n2854 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/la0/la_window_depth[3] ), 
            .O(\edb_top_inst/n2872 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4518 .LUTMASK = 16'hf305;
    EFX_LUT4 \edb_top_inst/LUT__4519  (.I0(\edb_top_inst/n2857 ), .I1(\edb_top_inst/la0/la_window_depth[2] ), 
            .I2(\edb_top_inst/la0/la_window_depth[4] ), .I3(\edb_top_inst/n2872 ), 
            .O(\edb_top_inst/n2873 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4519 .LUTMASK = 16'h000b;
    EFX_LUT4 \edb_top_inst/LUT__4520  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I2(\edb_top_inst/n2678 ), .I3(\edb_top_inst/n2873 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4520 .LUTMASK = 16'hff80;
    EFX_LUT4 \edb_top_inst/LUT__4521  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), .I2(\edb_top_inst/la0/la_window_depth[1] ), 
            .O(\edb_top_inst/n2874 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4521 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4522  (.I0(\edb_top_inst/n2874 ), .I1(\edb_top_inst/n2870 ), 
            .I2(\edb_top_inst/la0/la_window_depth[0] ), .O(\edb_top_inst/n2875 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4522 .LUTMASK = 16'hcaca;
    EFX_LUT4 \edb_top_inst/LUT__4523  (.I0(\edb_top_inst/n2875 ), .I1(\edb_top_inst/n2861 ), 
            .I2(\edb_top_inst/la0/la_window_depth[2] ), .I3(\edb_top_inst/n2690 ), 
            .O(\edb_top_inst/n2876 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4523 .LUTMASK = 16'hca00;
    EFX_LUT4 \edb_top_inst/LUT__4524  (.I0(\edb_top_inst/n2844 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/n2876 ), .O(\edb_top_inst/n2877 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4524 .LUTMASK = 16'h0b0b;
    EFX_LUT4 \edb_top_inst/LUT__4525  (.I0(\edb_top_inst/n2679 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] ), 
            .I2(\edb_top_inst/n2877 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_write_addr/out_phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f8f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4525 .LUTMASK = 16'h8f8f;
    EFX_LUT4 \edb_top_inst/LUT__4526  (.I0(\edb_top_inst/n2700 ), .I1(\edb_top_inst/n2838 ), 
            .I2(\edb_top_inst/n2837 ), .I3(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4526 .LUTMASK = 16'h8f88;
    EFX_LUT4 \edb_top_inst/LUT__4527  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I1(\edb_top_inst/n2839 ), .I2(\edb_top_inst/n2841 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4527 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4528  (.I0(\edb_top_inst/n2844 ), .I1(\edb_top_inst/n2700 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .I3(\edb_top_inst/n2842 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4528 .LUTMASK = 16'hf444;
    EFX_LUT4 \edb_top_inst/LUT__4529  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I1(\edb_top_inst/n2845 ), .I2(\edb_top_inst/n2848 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4529 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4530  (.I0(\edb_top_inst/n2850 ), .I1(\edb_top_inst/n2845 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I3(\edb_top_inst/n2853 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4530 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4531  (.I0(\edb_top_inst/n2849 ), .I1(\edb_top_inst/n2845 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I3(\edb_top_inst/n2858 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4531 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4532  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I1(\edb_top_inst/n2859 ), .I2(\edb_top_inst/n2862 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4532 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4533  (.I0(\edb_top_inst/n2678 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I2(\edb_top_inst/n2865 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8f8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4533 .LUTMASK = 16'hf8f8;
    EFX_LUT4 \edb_top_inst/LUT__4534  (.I0(\edb_top_inst/n2708 ), .I1(\edb_top_inst/n2678 ), 
            .I2(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I3(\edb_top_inst/n2869 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4534 .LUTMASK = 16'hff40;
    EFX_LUT4 \edb_top_inst/LUT__4535  (.I0(\edb_top_inst/la0/la_window_depth[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I2(\edb_top_inst/n2678 ), .I3(\edb_top_inst/n2873 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff80, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4535 .LUTMASK = 16'hff80;
    EFX_LUT4 \edb_top_inst/LUT__4536  (.I0(\edb_top_inst/n2679 ), .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] ), 
            .I2(\edb_top_inst/n2877 ), .O(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/transcode_read_addr/out_phy_addr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f8f, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4536 .LUTMASK = 16'h8f8f;
    EFX_LUT4 \edb_top_inst/LUT__4537  (.I0(\edb_top_inst/la0/module_state[1] ), 
            .I1(\edb_top_inst/la0/module_state[0] ), .I2(\edb_top_inst/la0/module_state[2] ), 
            .I3(\edb_top_inst/la0/module_state[3] ), .O(\edb_top_inst/n2878 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fb8, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4537 .LUTMASK = 16'h0fb8;
    EFX_LUT4 \edb_top_inst/LUT__4538  (.I0(\edb_top_inst/n2878 ), .I1(jtag_inst1_UPDATE), 
            .I2(\edb_top_inst/edb_user_dr[81] ), .I3(jtag_inst1_SEL), .O(\edb_top_inst/debug_hub_inst/n266 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4538 .LUTMASK = 16'h4000;
    EFX_LUT4 \edb_top_inst/LUT__4539  (.I0(jtag_inst1_SEL), .I1(jtag_inst1_SHIFT), 
            .O(\edb_top_inst/debug_hub_inst/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4539 .LUTMASK = 16'h8888;
    EFX_LUT4 \edb_top_inst/LUT__4540  (.I0(\edb_top_inst/la0/opcode[0] ), 
            .I1(\edb_top_inst/la0/opcode[3] ), .I2(\edb_top_inst/la0/opcode[2] ), 
            .I3(\edb_top_inst/la0/opcode[1] ), .O(\edb_top_inst/n2250 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000, EFX_ATTRIBUTE_INSTANCE__IS_STF_LUT=TRUE */ ;
    defparam \edb_top_inst/LUT__4540 .LUTMASK = 16'h1000;
    EFX_ADD \edb_top_inst/la0/add_91/i1  (.I0(\edb_top_inst/la0/address_counter[0] ), 
            .I1(\edb_top_inst/n1285 ), .CI(1'b0), .O(\edb_top_inst/n53 ), 
            .CO(\edb_top_inst/n54 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i1 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i2  (.I0(\edb_top_inst/la0/bit_count[1] ), 
            .I1(\edb_top_inst/la0/bit_count[0] ), .CI(1'b0), .O(\edb_top_inst/n55 ), 
            .CO(\edb_top_inst/n56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3689)
    defparam \edb_top_inst/la0/add_100/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[0] ), .CI(1'b0), 
            .O(\edb_top_inst/n341 ), .CO(\edb_top_inst/n342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4611)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/n774 ), .CO(\edb_top_inst/n775 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4618)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[0] ), 
            .CI(1'b0), .O(\edb_top_inst/n776 ), .CO(\edb_top_inst/n777 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4622)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[1] ), 
            .I1(\edb_top_inst/la0/la_biu_inst/fifo_counter[0] ), .CI(1'b0), 
            .O(\edb_top_inst/n778 ), .CO(\edb_top_inst/n779 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4629)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2  (.I0(\edb_top_inst/la0/la_sample_cnt[1] ), 
            .I1(\edb_top_inst/la0/la_sample_cnt[0] ), .CI(1'b0), .O(\edb_top_inst/n780 ), 
            .CO(\edb_top_inst/n781 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12  (.I0(\edb_top_inst/la0/la_sample_cnt[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n941 ), .O(\edb_top_inst/n939 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11  (.I0(\edb_top_inst/la0/la_sample_cnt[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n943 ), .O(\edb_top_inst/n940 ), 
            .CO(\edb_top_inst/n941 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10  (.I0(\edb_top_inst/la0/la_sample_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n945 ), .O(\edb_top_inst/n942 ), 
            .CO(\edb_top_inst/n943 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9  (.I0(\edb_top_inst/la0/la_sample_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n947 ), .O(\edb_top_inst/n944 ), 
            .CO(\edb_top_inst/n945 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8  (.I0(\edb_top_inst/la0/la_sample_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n949 ), .O(\edb_top_inst/n946 ), 
            .CO(\edb_top_inst/n947 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7  (.I0(\edb_top_inst/la0/la_sample_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n951 ), .O(\edb_top_inst/n948 ), 
            .CO(\edb_top_inst/n949 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6  (.I0(\edb_top_inst/la0/la_sample_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n953 ), .O(\edb_top_inst/n950 ), 
            .CO(\edb_top_inst/n951 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5  (.I0(\edb_top_inst/la0/la_sample_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n955 ), .O(\edb_top_inst/n952 ), 
            .CO(\edb_top_inst/n953 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4  (.I0(\edb_top_inst/la0/la_sample_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n957 ), .O(\edb_top_inst/n954 ), 
            .CO(\edb_top_inst/n955 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3  (.I0(\edb_top_inst/la0/la_sample_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n781 ), .O(\edb_top_inst/n956 ), 
            .CO(\edb_top_inst/n957 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4643)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_46/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/counter[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n960 ), .O(\edb_top_inst/n958 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4629)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n962 ), .O(\edb_top_inst/n959 ), 
            .CO(\edb_top_inst/n960 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4629)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n964 ), .O(\edb_top_inst/n961 ), 
            .CO(\edb_top_inst/n962 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4629)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n966 ), .O(\edb_top_inst/n963 ), 
            .CO(\edb_top_inst/n964 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4629)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n968 ), .O(\edb_top_inst/n965 ), 
            .CO(\edb_top_inst/n966 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4629)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n970 ), .O(\edb_top_inst/n967 ), 
            .CO(\edb_top_inst/n968 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4629)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n972 ), .O(\edb_top_inst/n969 ), 
            .CO(\edb_top_inst/n970 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4629)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n974 ), .O(\edb_top_inst/n971 ), 
            .CO(\edb_top_inst/n972 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4629)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n976 ), .O(\edb_top_inst/n973 ), 
            .CO(\edb_top_inst/n974 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4629)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_counter[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n779 ), .O(\edb_top_inst/n975 ), 
            .CO(\edb_top_inst/n976 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4629)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_21/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1002 ), .O(\edb_top_inst/n999 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4622)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1004 ), .O(\edb_top_inst/n1001 ), 
            .CO(\edb_top_inst/n1002 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4622)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1006 ), .O(\edb_top_inst/n1003 ), 
            .CO(\edb_top_inst/n1004 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4622)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1008 ), .O(\edb_top_inst/n1005 ), 
            .CO(\edb_top_inst/n1006 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4622)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1010 ), .O(\edb_top_inst/n1007 ), 
            .CO(\edb_top_inst/n1008 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4622)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1012 ), .O(\edb_top_inst/n1009 ), 
            .CO(\edb_top_inst/n1010 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4622)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1014 ), .O(\edb_top_inst/n1011 ), 
            .CO(\edb_top_inst/n1012 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4622)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1016 ), .O(\edb_top_inst/n1013 ), 
            .CO(\edb_top_inst/n1014 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4622)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_wr_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n777 ), .O(\edb_top_inst/n1015 ), 
            .CO(\edb_top_inst/n1016 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4622)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_12/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1051 ), .O(\edb_top_inst/n1048 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4618)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1053 ), .O(\edb_top_inst/n1050 ), 
            .CO(\edb_top_inst/n1051 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4618)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1055 ), .O(\edb_top_inst/n1052 ), 
            .CO(\edb_top_inst/n1053 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4618)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1057 ), .O(\edb_top_inst/n1054 ), 
            .CO(\edb_top_inst/n1055 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4618)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1059 ), .O(\edb_top_inst/n1056 ), 
            .CO(\edb_top_inst/n1057 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4618)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1061 ), .O(\edb_top_inst/n1058 ), 
            .CO(\edb_top_inst/n1059 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4618)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1063 ), .O(\edb_top_inst/n1060 ), 
            .CO(\edb_top_inst/n1061 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4618)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1065 ), .O(\edb_top_inst/n1062 ), 
            .CO(\edb_top_inst/n1063 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4618)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3  (.I0(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/segment_rd_pointer[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n775 ), .O(\edb_top_inst/n1064 ), 
            .CO(\edb_top_inst/n1065 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4618)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_10/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1068 ), .O(\edb_top_inst/n1066 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4611)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1070 ), .O(\edb_top_inst/n1067 ), 
            .CO(\edb_top_inst/n1068 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4611)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1072 ), .O(\edb_top_inst/n1069 ), 
            .CO(\edb_top_inst/n1070 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4611)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1074 ), .O(\edb_top_inst/n1071 ), 
            .CO(\edb_top_inst/n1072 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4611)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1076 ), .O(\edb_top_inst/n1073 ), 
            .CO(\edb_top_inst/n1074 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4611)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1078 ), .O(\edb_top_inst/n1075 ), 
            .CO(\edb_top_inst/n1076 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4611)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1080 ), .O(\edb_top_inst/n1077 ), 
            .CO(\edb_top_inst/n1078 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4611)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1082 ), .O(\edb_top_inst/n1079 ), 
            .CO(\edb_top_inst/n1080 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4611)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3  (.I0(\edb_top_inst/la0/la_biu_inst/la_window_fill_cnt[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n342 ), .O(\edb_top_inst/n1081 ), 
            .CO(\edb_top_inst/n1082 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(4611)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/add_9/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i6  (.I0(\edb_top_inst/la0/bit_count[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1085 ), .O(\edb_top_inst/n1083 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3689)
    defparam \edb_top_inst/la0/add_100/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i5  (.I0(\edb_top_inst/la0/bit_count[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1087 ), .O(\edb_top_inst/n1084 ), 
            .CO(\edb_top_inst/n1085 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3689)
    defparam \edb_top_inst/la0/add_100/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i4  (.I0(\edb_top_inst/la0/bit_count[3] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1089 ), .O(\edb_top_inst/n1086 ), 
            .CO(\edb_top_inst/n1087 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3689)
    defparam \edb_top_inst/la0/add_100/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_100/i3  (.I0(\edb_top_inst/la0/bit_count[2] ), 
            .I1(1'b0), .CI(\edb_top_inst/n56 ), .O(\edb_top_inst/n1088 ), 
            .CO(\edb_top_inst/n1089 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3689)
    defparam \edb_top_inst/la0/add_100/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_100/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i26  (.I0(\edb_top_inst/la0/address_counter[25] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1104 ), .O(\edb_top_inst/n1101 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i26 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i25  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1106 ), .O(\edb_top_inst/n1103 ), 
            .CO(\edb_top_inst/n1104 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i25 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i24  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1108 ), .O(\edb_top_inst/n1105 ), 
            .CO(\edb_top_inst/n1106 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i24 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i23  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1110 ), .O(\edb_top_inst/n1107 ), 
            .CO(\edb_top_inst/n1108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i23 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i22  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1112 ), .O(\edb_top_inst/n1109 ), 
            .CO(\edb_top_inst/n1110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i22 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i21  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1114 ), .O(\edb_top_inst/n1111 ), 
            .CO(\edb_top_inst/n1112 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i21 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i20  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1116 ), .O(\edb_top_inst/n1113 ), 
            .CO(\edb_top_inst/n1114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i20 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i19  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1118 ), .O(\edb_top_inst/n1115 ), 
            .CO(\edb_top_inst/n1116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i19 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i18  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1120 ), .O(\edb_top_inst/n1117 ), 
            .CO(\edb_top_inst/n1118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i18 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i17  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1122 ), .O(\edb_top_inst/n1119 ), 
            .CO(\edb_top_inst/n1120 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i17 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i16  (.I0(\edb_top_inst/la0/address_counter[15] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1124 ), .O(\edb_top_inst/n1121 ), 
            .CO(\edb_top_inst/n1122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i16 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i15  (.I0(\edb_top_inst/la0/address_counter[14] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1126 ), .O(\edb_top_inst/n1123 ), 
            .CO(\edb_top_inst/n1124 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i15 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i14  (.I0(\edb_top_inst/la0/address_counter[13] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1128 ), .O(\edb_top_inst/n1125 ), 
            .CO(\edb_top_inst/n1126 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i14 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i13  (.I0(\edb_top_inst/la0/address_counter[12] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1130 ), .O(\edb_top_inst/n1127 ), 
            .CO(\edb_top_inst/n1128 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i13 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i12  (.I0(\edb_top_inst/la0/address_counter[11] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1132 ), .O(\edb_top_inst/n1129 ), 
            .CO(\edb_top_inst/n1130 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i12 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i11  (.I0(\edb_top_inst/la0/address_counter[10] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1134 ), .O(\edb_top_inst/n1131 ), 
            .CO(\edb_top_inst/n1132 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i10  (.I0(\edb_top_inst/la0/address_counter[9] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1136 ), .O(\edb_top_inst/n1133 ), 
            .CO(\edb_top_inst/n1134 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i9  (.I0(\edb_top_inst/la0/address_counter[8] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1138 ), .O(\edb_top_inst/n1135 ), 
            .CO(\edb_top_inst/n1136 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i8  (.I0(\edb_top_inst/la0/address_counter[7] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1140 ), .O(\edb_top_inst/n1137 ), 
            .CO(\edb_top_inst/n1138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i7  (.I0(\edb_top_inst/la0/address_counter[6] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1142 ), .O(\edb_top_inst/n1139 ), 
            .CO(\edb_top_inst/n1140 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i6  (.I0(\edb_top_inst/la0/address_counter[5] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1144 ), .O(\edb_top_inst/n1141 ), 
            .CO(\edb_top_inst/n1142 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i5  (.I0(\edb_top_inst/la0/address_counter[4] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1146 ), .O(\edb_top_inst/n1143 ), 
            .CO(\edb_top_inst/n1144 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i4  (.I0(\edb_top_inst/la0/address_counter[3] ), 
            .I1(\edb_top_inst/n2244 ), .CI(\edb_top_inst/n1148 ), .O(\edb_top_inst/n1145 ), 
            .CO(\edb_top_inst/n1146 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i3  (.I0(\edb_top_inst/la0/address_counter[2] ), 
            .I1(\edb_top_inst/n2247 ), .CI(\edb_top_inst/n1150 ), .O(\edb_top_inst/n1147 ), 
            .CO(\edb_top_inst/n1148 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_91/i2  (.I0(\edb_top_inst/la0/address_counter[1] ), 
            .I1(\edb_top_inst/n2250 ), .CI(\edb_top_inst/n54 ), .O(\edb_top_inst/n1149 ), 
            .CO(\edb_top_inst/n1150 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3662)
    defparam \edb_top_inst/la0/add_91/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_91/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i11  (.I0(\edb_top_inst/la0/address_counter[25] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1165 ), .O(\edb_top_inst/n1162 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3661)
    defparam \edb_top_inst/la0/add_90/i11 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i10  (.I0(\edb_top_inst/la0/address_counter[24] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1167 ), .O(\edb_top_inst/n1164 ), 
            .CO(\edb_top_inst/n1165 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3661)
    defparam \edb_top_inst/la0/add_90/i10 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i9  (.I0(\edb_top_inst/la0/address_counter[23] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1169 ), .O(\edb_top_inst/n1166 ), 
            .CO(\edb_top_inst/n1167 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3661)
    defparam \edb_top_inst/la0/add_90/i9 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i8  (.I0(\edb_top_inst/la0/address_counter[22] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1171 ), .O(\edb_top_inst/n1168 ), 
            .CO(\edb_top_inst/n1169 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3661)
    defparam \edb_top_inst/la0/add_90/i8 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i7  (.I0(\edb_top_inst/la0/address_counter[21] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1173 ), .O(\edb_top_inst/n1170 ), 
            .CO(\edb_top_inst/n1171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3661)
    defparam \edb_top_inst/la0/add_90/i7 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i6  (.I0(\edb_top_inst/la0/address_counter[20] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1178 ), .O(\edb_top_inst/n1172 ), 
            .CO(\edb_top_inst/n1173 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3661)
    defparam \edb_top_inst/la0/add_90/i6 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i5  (.I0(\edb_top_inst/la0/address_counter[19] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1180 ), .O(\edb_top_inst/n1177 ), 
            .CO(\edb_top_inst/n1178 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3661)
    defparam \edb_top_inst/la0/add_90/i5 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i4  (.I0(\edb_top_inst/la0/address_counter[18] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1182 ), .O(\edb_top_inst/n1179 ), 
            .CO(\edb_top_inst/n1180 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3661)
    defparam \edb_top_inst/la0/add_90/i4 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i3  (.I0(\edb_top_inst/la0/address_counter[17] ), 
            .I1(1'b0), .CI(\edb_top_inst/n1184 ), .O(\edb_top_inst/n1181 ), 
            .CO(\edb_top_inst/n1182 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3661)
    defparam \edb_top_inst/la0/add_90/i3 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \edb_top_inst/la0/add_90/i2  (.I0(\edb_top_inst/la0/address_counter[16] ), 
            .I1(\edb_top_inst/la0/address_counter[15] ), .CI(1'b0), .O(\edb_top_inst/n1183 ), 
            .CO(\edb_top_inst/n1184 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_ADD=TRUE */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(3661)
    defparam \edb_top_inst/la0/add_90/i2 .I0_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/add_90/i2 .I1_POLARITY = 1'b1;
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[0] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[1] , \edb_top_inst/la0/la_biu_inst/fifo_dout[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=df1292e9 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[2] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[3] , \edb_top_inst/la0/la_biu_inst/fifo_dout[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=d7b17582 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[4] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[5] , \edb_top_inst/la0/la_biu_inst/fifo_dout[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=3eae9e73 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[6] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[7] , \edb_top_inst/la0/la_biu_inst/fifo_dout[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=80ce81b6 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[8] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[9] , \edb_top_inst/la0/la_biu_inst/fifo_dout[8] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=68cb4782 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[11] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[10] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[11] , \edb_top_inst/la0/la_biu_inst/fifo_dout[10] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=0105c037 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[13] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[12] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[13] , \edb_top_inst/la0/la_biu_inst/fifo_dout[12] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=a9e573bd */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[15] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[14] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[15] , \edb_top_inst/la0/la_biu_inst/fifo_dout[14] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=d5089fa5 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$g12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[17] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[16] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[17] , \edb_top_inst/la0/la_biu_inst/fifo_dout[16] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=f5556ccb */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$h12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[19] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[18] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[19] , \edb_top_inst/la0/la_biu_inst/fifo_dout[18] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=7dedc663 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$i12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[21] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[20] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[21] , \edb_top_inst/la0/la_biu_inst/fifo_dout[20] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=128f5a70 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$j12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[23] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[22] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[23] , \edb_top_inst/la0/la_biu_inst/fifo_dout[22] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=d8939b8d */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$k12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[25] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[24] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[25] , \edb_top_inst/la0/la_biu_inst/fifo_dout[24] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=63be41e7 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$l12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[27] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[26] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[27] , \edb_top_inst/la0/la_biu_inst/fifo_dout[26] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=b6f477c9 */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$m12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1  (.WCLK(\clk~O ), 
            .RCLK(\clk~O ), .WCLKE(1'b1), .WE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/push_p2 ), 
            .RE(\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/n658 ), 
            .WDATA({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[29] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/din_p2[28] }), 
            .WADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/wr_pointer[0] }), 
            .RADDR({\edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[10] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[9] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[8] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[7] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[6] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[5] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[4] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[3] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[2] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[1] , 
            \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/phy_addr[0] }), 
            .RDATA({\edb_top_inst/la0/la_biu_inst/fifo_dout[29] , \edb_top_inst/la0/la_biu_inst/fifo_dout[28] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b1, EFX_ATTRIBUTE_INSTANCE__IS_STF_RAM_5K=TRUE, EFX_ATTRIBUTE_NET__RAMINFO_ID=ef93be5b */ ;   // /home/amritansh/Downloads/efinity/2023.1/project/Dual_TX_Controller/work_dbg/debug_top.v(418)
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .READ_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .WRITE_WIDTH = 2;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .WCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .WCLKE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .WE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .RCLK_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .RE_POLARITY = 1'b1;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .OUTPUT_REG = 1'b0;
    defparam \edb_top_inst/la0/la_biu_inst/fifo_with_read_inst/simple_dual_port_ram_inst/ram__D$n1 .WRITE_MODE = "READ_FIRST";
    EFX_LUT4 LUT__6746 (.I0(ceg_net133), .I1(\state[0] ), .O(ceg_net108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__6746.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__6747 (.I0(\i[1] ), .I1(\i[0] ), .I2(\data_length[1] ), 
            .I3(\data_length[0] ), .O(n4503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__6747.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__6748 (.I0(\data_length[4] ), .I1(\i[4] ), .I2(\data_length[3] ), 
            .I3(\i[3] ), .O(n4504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__6748.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__6749 (.I0(\i[2] ), .I1(n4503), .I2(\data_length[2] ), 
            .I3(n4504), .O(n4505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7100 */ ;
    defparam LUT__6749.LUTMASK = 16'h7100;
    EFX_LUT4 LUT__6750 (.I0(\i[4] ), .I1(\i[3] ), .I2(\data_length[4] ), 
            .I3(\data_length[3] ), .O(n4506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8eaf */ ;
    defparam LUT__6750.LUTMASK = 16'h8eaf;
    EFX_LUT4 LUT__6751 (.I0(\i[5] ), .I1(\data_length[5] ), .I2(n4505), 
            .I3(n4506), .O(n4507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4dd */ ;
    defparam LUT__6751.LUTMASK = 16'hd4dd;
    EFX_LUT4 LUT__6752 (.I0(ceg_net108), .I1(n4507), .O(ceg_net98)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__6752.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__6753 (.I0(ceg_net133), .I1(n4507), .I2(\state[1] ), 
            .I3(\state[0] ), .O(ceg_net127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbb0f */ ;
    defparam LUT__6753.LUTMASK = 16'hbb0f;
    EFX_LUT4 LUT__6754 (.I0(n4507), .I1(\state[0] ), .I2(ceg_net133), 
            .O(ceg_net130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__6754.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__6755 (.I0(\state[0] ), .I1(n4507), .O(n257_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6755.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6756 (.I0(\i[0] ), .I1(n4507), .O(n62_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6756.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6757 (.I0(RX_DV), .I1(\uart_rx/r_RX_Byte[6] ), .O(\received_data[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6757.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6758 (.I0(RX_DV), .I1(\uart_rx/r_RX_Byte[7] ), .O(\received_data[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6758.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6759 (.I0(\received_data[6] ), .I1(\received_data[7] ), 
            .O(\equal_4/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__6759.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__6760 (.I0(\state[0] ), .I1(ceg_net133), .O(ceg_net120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__6760.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__6761 (.I0(RX_DV), .I1(\state[1] ), .O(ceg_net138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6761.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6762 (.I0(\uart_rx/r_Clock_Count[4] ), .I1(\uart_rx/r_Clock_Count[6] ), 
            .I2(\uart_rx/r_Clock_Count[5] ), .I3(\uart_rx/r_Clock_Count[3] ), 
            .O(n4508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6762.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6763 (.I0(\uart_rx/r_Clock_Count[0] ), .I1(\uart_rx/r_Clock_Count[1] ), 
            .O(n4509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6763.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6764 (.I0(\uart_rx/r_Clock_Count[2] ), .I1(\uart_rx/r_Clock_Count[7] ), 
            .I2(n4508), .I3(n4509), .O(n4510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6764.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6765 (.I0(\uart_rx/r_Clock_Count[2] ), .I1(\uart_rx/r_Clock_Count[1] ), 
            .I2(\uart_rx/r_Clock_Count[3] ), .I3(\uart_rx/r_Clock_Count[4] ), 
            .O(n4511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6765.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6766 (.I0(\uart_rx/r_Clock_Count[5] ), .I1(n4511), .I2(\uart_rx/r_Clock_Count[6] ), 
            .I3(\uart_rx/r_Clock_Count[7] ), .O(\uart_rx/n43 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__6766.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__6767 (.I0(n4510), .I1(\uart_rx/r_SM_Main[0] ), .I2(\uart_rx/n43 ), 
            .I3(\uart_rx/r_SM_Main[1] ), .O(n4512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__6767.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__6768 (.I0(\uart_rx/r_Clock_Count[0] ), .I1(n4512), .O(\uart_rx/n375 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6768.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6769 (.I0(rx), .I1(\uart_rx/r_SM_Main[0] ), .O(n4513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6769.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6770 (.I0(\uart_rx/r_SM_Main[1] ), .I1(n4510), .I2(n4513), 
            .I3(\uart_rx/r_SM_Main[2] ), .O(ceg_net78)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff40 */ ;
    defparam LUT__6770.LUTMASK = 16'hff40;
    EFX_LUT4 LUT__6771 (.I0(\uart_rx/r_SM_Main[2] ), .I1(\uart_rx/r_SM_Main[1] ), 
            .O(\uart_rx/n407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6771.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6772 (.I0(\uart_rx/r_SM_Main[2] ), .I1(\uart_rx/n43 ), 
            .I2(\uart_rx/r_SM_Main[0] ), .I3(\uart_rx/r_SM_Main[1] ), .O(ceg_net153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heff0 */ ;
    defparam LUT__6772.LUTMASK = 16'heff0;
    EFX_LUT4 LUT__6773 (.I0(\uart_rx/r_Bit_Index[0] ), .I1(\uart_rx/r_Bit_Index[1] ), 
            .I2(\uart_rx/r_Bit_Index[2] ), .I3(\uart_rx/r_SM_Main[1] ), 
            .O(n4514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6773.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6774 (.I0(\uart_rx/r_SM_Main[0] ), .I1(\uart_rx/n43 ), 
            .I2(n4514), .O(\uart_rx/n444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6774.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6775 (.I0(\uart_rx/r_Bit_Index[0] ), .I1(\uart_rx/r_SM_Main[1] ), 
            .O(\uart_rx/n382 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6775.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6776 (.I0(\uart_rx/n43 ), .I1(\uart_rx/r_SM_Main[1] ), 
            .I2(\uart_rx/r_SM_Main[2] ), .I3(\uart_rx/r_SM_Main[0] ), .O(ceg_net146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__6776.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__6777 (.I0(\uart_rx/r_Bit_Index[0] ), .I1(\uart_rx/r_Bit_Index[1] ), 
            .I2(\uart_rx/r_Bit_Index[2] ), .O(n4515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6777.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6778 (.I0(\uart_rx/n43 ), .I1(n4515), .I2(rx), .I3(\uart_rx/r_SM_Main[1] ), 
            .O(n4516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__6778.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__6779 (.I0(n4516), .I1(n4512), .I2(\uart_rx/r_SM_Main[0] ), 
            .O(\uart_rx/n372 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6779.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6780 (.I0(n4512), .I1(\uart_rx/r_Clock_Count[0] ), .I2(\uart_rx/r_Clock_Count[1] ), 
            .O(\uart_rx/n316 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__6780.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__6781 (.I0(n4512), .I1(\uart_rx/r_Clock_Count[2] ), .I2(n4509), 
            .O(\uart_rx/n319 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__6781.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__6782 (.I0(\uart_rx/r_Clock_Count[2] ), .I1(n4509), .I2(n4512), 
            .I3(\uart_rx/r_Clock_Count[3] ), .O(\uart_rx/n322 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__6782.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__6783 (.I0(\uart_rx/r_Clock_Count[2] ), .I1(\uart_rx/r_Clock_Count[3] ), 
            .I2(n4509), .O(n4517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6783.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6784 (.I0(n4512), .I1(\uart_rx/r_Clock_Count[4] ), .I2(n4517), 
            .O(\uart_rx/n325 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__6784.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__6785 (.I0(\uart_rx/r_Clock_Count[4] ), .I1(n4517), .I2(n4512), 
            .I3(\uart_rx/r_Clock_Count[5] ), .O(\uart_rx/n328 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__6785.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__6786 (.I0(\uart_rx/r_Clock_Count[4] ), .I1(\uart_rx/r_Clock_Count[5] ), 
            .I2(n4517), .O(n4518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6786.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6787 (.I0(n4512), .I1(\uart_rx/r_Clock_Count[6] ), .I2(n4518), 
            .O(\uart_rx/n331 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__6787.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__6788 (.I0(\uart_rx/r_Clock_Count[6] ), .I1(n4518), .I2(n4512), 
            .I3(\uart_rx/r_Clock_Count[7] ), .O(\uart_rx/n334 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__6788.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__6789 (.I0(\uart_rx/r_SM_Main[0] ), .I1(\uart_rx/n43 ), 
            .I2(\uart_rx/n407 ), .O(n4519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6789.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6790 (.I0(\uart_rx/r_Bit_Index[1] ), .I1(\uart_rx/r_Bit_Index[2] ), 
            .I2(\uart_rx/r_Bit_Index[0] ), .I3(n4519), .O(\uart_rx/n429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6790.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6791 (.I0(\uart_rx/r_Bit_Index[0] ), .I1(\uart_rx/r_Bit_Index[2] ), 
            .I2(\uart_rx/r_Bit_Index[1] ), .I3(n4519), .O(\uart_rx/n431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6791.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6792 (.I0(\uart_rx/r_Bit_Index[2] ), .I1(\uart_rx/r_Bit_Index[1] ), 
            .I2(\uart_rx/r_Bit_Index[0] ), .I3(n4519), .O(\uart_rx/n433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6792.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6793 (.I0(\uart_rx/r_Bit_Index[0] ), .I1(\uart_rx/r_Bit_Index[1] ), 
            .I2(\uart_rx/r_Bit_Index[2] ), .I3(n4519), .O(\uart_rx/n435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6793.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6794 (.I0(\uart_rx/r_Bit_Index[1] ), .I1(\uart_rx/r_Bit_Index[0] ), 
            .I2(\uart_rx/r_Bit_Index[2] ), .I3(n4519), .O(\uart_rx/n437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6794.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6795 (.I0(\uart_rx/r_Bit_Index[0] ), .I1(\uart_rx/r_Bit_Index[1] ), 
            .I2(\uart_rx/r_Bit_Index[2] ), .I3(n4519), .O(\uart_rx/n439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6795.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6796 (.I0(n4515), .I1(n4519), .O(\uart_rx/n441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6796.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6797 (.I0(\uart_rx/r_Bit_Index[0] ), .I1(\uart_rx/r_Bit_Index[1] ), 
            .I2(\uart_rx/r_SM_Main[1] ), .O(\uart_rx/n359 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6797.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6798 (.I0(\uart_rx/r_Bit_Index[0] ), .I1(\uart_rx/r_Bit_Index[1] ), 
            .I2(\uart_rx/r_Bit_Index[2] ), .I3(\uart_rx/r_SM_Main[1] ), 
            .O(\uart_rx/n363 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__6798.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6799 (.I0(rx), .I1(\uart_rx/r_SM_Main[0] ), .I2(n4510), 
            .O(n4520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6799.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6800 (.I0(\uart_rx/n43 ), .I1(\uart_rx/r_SM_Main[0] ), 
            .I2(n4520), .I3(\uart_rx/r_SM_Main[1] ), .O(\uart_rx/n309 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__6800.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__6801 (.I0(\uart_rx/r_SM_Main[0] ), .I1(\uart_rx/r_SM_Main[1] ), 
            .O(\uart_rx/n385 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6801.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6802 (.I0(RX_DV), .I1(\uart_rx/r_RX_Byte[1] ), .O(\received_data[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6802.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6803 (.I0(RX_DV), .I1(\uart_rx/r_RX_Byte[2] ), .O(\received_data[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6803.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6804 (.I0(RX_DV), .I1(\uart_rx/r_RX_Byte[3] ), .O(\received_data[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6804.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6805 (.I0(RX_DV), .I1(\uart_rx/r_RX_Byte[4] ), .O(\received_data[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6805.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6806 (.I0(RX_DV), .I1(\uart_rx/r_RX_Byte[5] ), .O(\received_data[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6806.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6807 (.I0(\i[0] ), .I1(\i[1] ), .I2(n4507), .O(n61_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6807.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6808 (.I0(\i[0] ), .I1(\i[1] ), .O(n4521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6808.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6809 (.I0(\i[2] ), .I1(n4521), .I2(n4507), .O(n60_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6809.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6810 (.I0(\i[2] ), .I1(n4521), .I2(\i[3] ), .I3(n4507), 
            .O(n59_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__6810.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6811 (.I0(\i[2] ), .I1(\i[3] ), .I2(n4521), .O(n4522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6811.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6812 (.I0(\i[4] ), .I1(n4522), .I2(n4507), .O(n58_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6812.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6813 (.I0(\i[4] ), .I1(n4522), .I2(\i[5] ), .I3(n4507), 
            .O(n57)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__6813.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6814 (.I0(\uart_rx/r_RX_Byte[7] ), .I1(\received_data[6] ), 
            .O(\equal_5/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__6814.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__6815 (.I0(\uart_tx1/r_Clock_Count[2] ), .I1(\uart_tx1/r_Clock_Count[1] ), 
            .I2(\uart_tx1/r_Clock_Count[3] ), .I3(\uart_tx1/r_Clock_Count[4] ), 
            .O(n4523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6815.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6816 (.I0(n4523), .I1(\uart_tx1/r_Clock_Count[5] ), .I2(\uart_tx1/r_Clock_Count[6] ), 
            .O(n4524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6816.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6817 (.I0(\uart_tx1/r_SM_Main[1] ), .I1(\uart_tx1/r_SM_Main[0] ), 
            .I2(n4524), .O(n4525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__6817.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__6818 (.I0(\uart_tx1/r_Clock_Count[0] ), .I1(n4525), .O(\uart_tx1/n119 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6818.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6819 (.I0(\uart_tx1/r_TX_Data[7] ), .I1(\uart_tx1/r_TX_Data[5] ), 
            .I2(\uart_tx1/r_Bit_Index[0] ), .I3(\uart_tx1/r_Bit_Index[1] ), 
            .O(n4526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6819.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6820 (.I0(\uart_tx1/r_TX_Data[6] ), .I1(\uart_tx1/r_TX_Data[4] ), 
            .I2(\uart_tx1/r_Bit_Index[0] ), .I3(n4526), .O(n4527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6820.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6821 (.I0(\uart_tx1/r_TX_Data[3] ), .I1(\uart_tx1/r_TX_Data[1] ), 
            .I2(\uart_tx1/r_Bit_Index[0] ), .I3(\uart_tx1/r_Bit_Index[1] ), 
            .O(n4528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6821.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6822 (.I0(\uart_tx1/r_TX_Data[2] ), .I1(\uart_tx1/r_TX_Data[0] ), 
            .I2(\uart_tx1/r_Bit_Index[0] ), .I3(n4528), .O(n4529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6822.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6823 (.I0(n4529), .I1(n4527), .I2(\uart_tx1/r_Bit_Index[2] ), 
            .O(n4530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6823.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6824 (.I0(n4530), .I1(\uart_tx1/r_SM_Main[0] ), .I2(\uart_tx1/r_SM_Main[1] ), 
            .O(\uart_tx1/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__6824.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__6825 (.I0(\uart_tx1/r_SM_Main[0] ), .I1(\uart_tx1/r_Bit_Index[0] ), 
            .I2(n4524), .I3(\uart_tx1/r_SM_Main[1] ), .O(\uart_tx1/select_38/Select_0/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400 */ ;
    defparam LUT__6825.LUTMASK = 16'h1400;
    EFX_LUT4 LUT__6827 (.I0(\uart_tx1/r_SM_Main[0] ), .I1(\uart_tx1/r_SM_Main[1] ), 
            .I2(DV), .O(\uart_tx1/n338 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6827.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6829 (.I0(\transmitter_select[1] ), .I1(\transmitter_select[0] ), 
            .O(n4532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6829.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6830 (.I0(\data[0] ), .I1(n4532), .O(\data_to_transmitter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6830.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6831 (.I0(n4523), .I1(\uart_tx1/r_Clock_Count[5] ), .I2(\uart_tx1/r_Clock_Count[6] ), 
            .I3(\uart_tx1/r_Bit_Index[0] ), .O(n4533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__6831.LUTMASK = 16'he000;
    EFX_LUT4 LUT__6832 (.I0(\uart_tx1/r_Bit_Index[1] ), .I1(\uart_tx1/r_Bit_Index[2] ), 
            .I2(\uart_tx1/r_SM_Main[1] ), .I3(n4533), .O(n4534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6832.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6833 (.I0(\uart_tx1/n338 ), .I1(n4534), .I2(n4524), 
            .I3(\uart_tx1/r_SM_Main[0] ), .O(\uart_tx1/n138 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__6833.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__6834 (.I0(\uart_tx1/r_Clock_Count[0] ), .I1(\uart_tx1/r_Clock_Count[1] ), 
            .I2(n4525), .O(\uart_tx1/n118 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6834.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6835 (.I0(\uart_tx1/r_Clock_Count[0] ), .I1(\uart_tx1/r_Clock_Count[1] ), 
            .O(n4535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6835.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6836 (.I0(\uart_tx1/r_Clock_Count[2] ), .I1(n4535), .I2(n4525), 
            .O(\uart_tx1/n117 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6836.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6837 (.I0(\uart_tx1/r_Clock_Count[2] ), .I1(n4535), .I2(\uart_tx1/r_Clock_Count[3] ), 
            .I3(n4525), .O(\uart_tx1/n116 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__6837.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6838 (.I0(\uart_tx1/r_Clock_Count[2] ), .I1(\uart_tx1/r_Clock_Count[3] ), 
            .I2(n4535), .O(n4536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6838.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6839 (.I0(\uart_tx1/r_Clock_Count[4] ), .I1(n4536), .I2(n4525), 
            .O(\uart_tx1/n115 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6839.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6840 (.I0(\uart_tx1/r_Clock_Count[4] ), .I1(n4536), .O(n4537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6840.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6841 (.I0(\uart_tx1/r_Clock_Count[5] ), .I1(n4537), .I2(n4525), 
            .O(\uart_tx1/n114 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6841.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6842 (.I0(\uart_tx1/r_Clock_Count[5] ), .I1(n4537), .I2(\uart_tx1/r_Clock_Count[6] ), 
            .I3(n4525), .O(\uart_tx1/n113 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6842.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6843 (.I0(\uart_tx1/r_SM_Main[0] ), .I1(n4533), .I2(\uart_tx1/r_SM_Main[1] ), 
            .I3(\uart_tx1/r_Bit_Index[1] ), .O(\uart_tx1/n122 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hba40 */ ;
    defparam LUT__6843.LUTMASK = 16'hba40;
    EFX_LUT4 LUT__6844 (.I0(\uart_tx1/r_Bit_Index[1] ), .I1(n4533), .O(n4538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6844.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6845 (.I0(\uart_tx1/r_SM_Main[0] ), .I1(n4538), .I2(\uart_tx1/r_SM_Main[1] ), 
            .I3(\uart_tx1/r_Bit_Index[2] ), .O(\uart_tx1/n121 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hba40 */ ;
    defparam LUT__6845.LUTMASK = 16'hba40;
    EFX_LUT4 LUT__6846 (.I0(\data[1] ), .I1(n4532), .O(\data_to_transmitter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6846.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6847 (.I0(\data[2] ), .I1(n4532), .O(\data_to_transmitter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6847.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6848 (.I0(\data[3] ), .I1(n4532), .O(\data_to_transmitter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6848.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6849 (.I0(\data[4] ), .I1(n4532), .O(\data_to_transmitter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6849.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6850 (.I0(\data[5] ), .I1(n4532), .O(\data_to_transmitter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6850.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6851 (.I0(\data[6] ), .I1(n4532), .O(\data_to_transmitter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6851.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6852 (.I0(\data[7] ), .I1(n4532), .O(\data_to_transmitter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6852.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6853 (.I0(\uart_tx1/r_SM_Main[0] ), .I1(n4524), .I2(\uart_tx1/r_SM_Main[1] ), 
            .O(\uart_tx1/n137 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__6853.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__6854 (.I0(\uart_tx2/r_TX_Data[7] ), .I1(\uart_tx2/r_TX_Data[5] ), 
            .I2(\uart_tx1/r_Bit_Index[0] ), .I3(\uart_tx1/r_Bit_Index[1] ), 
            .O(n4539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6854.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6855 (.I0(\uart_tx2/r_TX_Data[6] ), .I1(\uart_tx2/r_TX_Data[4] ), 
            .I2(\uart_tx1/r_Bit_Index[0] ), .I3(n4539), .O(n4540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6855.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6856 (.I0(\uart_tx2/r_TX_Data[3] ), .I1(\uart_tx2/r_TX_Data[1] ), 
            .I2(\uart_tx1/r_Bit_Index[0] ), .I3(\uart_tx1/r_Bit_Index[1] ), 
            .O(n4541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6856.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6857 (.I0(\uart_tx2/r_TX_Data[2] ), .I1(\uart_tx2/r_TX_Data[0] ), 
            .I2(\uart_tx1/r_Bit_Index[0] ), .I3(n4541), .O(n4542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6857.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6858 (.I0(n4542), .I1(n4540), .I2(\uart_tx1/r_Bit_Index[2] ), 
            .O(n4543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6858.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6859 (.I0(n4543), .I1(\uart_tx1/r_SM_Main[0] ), .I2(\uart_tx1/r_SM_Main[1] ), 
            .O(\uart_tx2/n110 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__6859.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__6860 (.I0(n4532), .I1(\data[0] ), .O(\data_to_transmitter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6860.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6861 (.I0(n4532), .I1(\data[1] ), .O(\data_to_transmitter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6861.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6862 (.I0(n4532), .I1(\data[2] ), .O(\data_to_transmitter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6862.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6863 (.I0(n4532), .I1(\data[3] ), .O(\data_to_transmitter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6863.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6864 (.I0(n4532), .I1(\data[4] ), .O(\data_to_transmitter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6864.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6865 (.I0(n4532), .I1(\data[5] ), .O(\data_to_transmitter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6865.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6866 (.I0(n4532), .I1(\data[6] ), .O(\data_to_transmitter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6866.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6867 (.I0(n4532), .I1(\data[7] ), .O(\data_to_transmitter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6867.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6744 (.I0(RX_DV), .I1(\uart_rx/r_RX_Byte[0] ), .O(\received_data[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6744.LUTMASK = 16'h8888;
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(clk), .O(\clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(jtag_inst1_TCK), .O(\jtag_inst1_TCK~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_f7a76cbb_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_f7a76cbb_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_f7a76cbb__2_2_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_f7a76cbb_185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_f7a76cbb_0
// module not written out since it is a black box. 
//

